library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity coeff_rom is
    generic(
        A_WIDTH : integer;
        D_WIDTH : integer
        );
    port (
        clk    : in  std_logic;
        clk_en : in  std_logic;
        addr   : in  unsigned(A_WIDTH - 1 downto 0);
        data   : out signed(D_WIDTH - 1 downto 0)
        );
end;

architecture rtl of coeff_rom is

    type t_coeff_list is array(0 to 2 ** A_WIDTH - 1) of
        signed(D_WIDTH - 1 downto 0);

    signal coeff_list : t_coeff_list := (
        to_signed(-144, D_WIDTH),
        to_signed(-142, D_WIDTH),
        to_signed(-140, D_WIDTH),
        to_signed(-138, D_WIDTH),
        to_signed(-136, D_WIDTH),
        to_signed(-134, D_WIDTH),
        to_signed(-132, D_WIDTH),
        to_signed(-129, D_WIDTH),
        to_signed(-127, D_WIDTH),
        to_signed(-125, D_WIDTH),
        to_signed(-122, D_WIDTH),
        to_signed(-120, D_WIDTH),
        to_signed(-117, D_WIDTH),
        to_signed(-115, D_WIDTH),
        to_signed(-112, D_WIDTH),
        to_signed(-110, D_WIDTH),
        to_signed(-107, D_WIDTH),
        to_signed(-104, D_WIDTH),
        to_signed(-102, D_WIDTH),
        to_signed(-99, D_WIDTH),
        to_signed(-96, D_WIDTH),
        to_signed(-93, D_WIDTH),
        to_signed(-90, D_WIDTH),
        to_signed(-87, D_WIDTH),
        to_signed(-84, D_WIDTH),
        to_signed(-81, D_WIDTH),
        to_signed(-78, D_WIDTH),
        to_signed(-75, D_WIDTH),
        to_signed(-72, D_WIDTH),
        to_signed(-69, D_WIDTH),
        to_signed(-66, D_WIDTH),
        to_signed(-63, D_WIDTH),
        to_signed(-59, D_WIDTH),
        to_signed(-56, D_WIDTH),
        to_signed(-53, D_WIDTH),
        to_signed(-50, D_WIDTH),
        to_signed(-46, D_WIDTH),
        to_signed(-43, D_WIDTH),
        to_signed(-40, D_WIDTH),
        to_signed(-36, D_WIDTH),
        to_signed(-33, D_WIDTH),
        to_signed(-29, D_WIDTH),
        to_signed(-26, D_WIDTH),
        to_signed(-22, D_WIDTH),
        to_signed(-19, D_WIDTH),
        to_signed(-15, D_WIDTH),
        to_signed(-12, D_WIDTH),
        to_signed(-8, D_WIDTH),
        to_signed(-5, D_WIDTH),
        to_signed(-1, D_WIDTH),
        to_signed(2, D_WIDTH),
        to_signed(6, D_WIDTH),
        to_signed(10, D_WIDTH),
        to_signed(13, D_WIDTH),
        to_signed(17, D_WIDTH),
        to_signed(20, D_WIDTH),
        to_signed(24, D_WIDTH),
        to_signed(28, D_WIDTH),
        to_signed(31, D_WIDTH),
        to_signed(35, D_WIDTH),
        to_signed(39, D_WIDTH),
        to_signed(42, D_WIDTH),
        to_signed(46, D_WIDTH),
        to_signed(49, D_WIDTH),
        to_signed(53, D_WIDTH),
        to_signed(57, D_WIDTH),
        to_signed(60, D_WIDTH),
        to_signed(64, D_WIDTH),
        to_signed(67, D_WIDTH),
        to_signed(71, D_WIDTH),
        to_signed(75, D_WIDTH),
        to_signed(78, D_WIDTH),
        to_signed(82, D_WIDTH),
        to_signed(85, D_WIDTH),
        to_signed(89, D_WIDTH),
        to_signed(92, D_WIDTH),
        to_signed(96, D_WIDTH),
        to_signed(99, D_WIDTH),
        to_signed(103, D_WIDTH),
        to_signed(106, D_WIDTH),
        to_signed(109, D_WIDTH),
        to_signed(113, D_WIDTH),
        to_signed(116, D_WIDTH),
        to_signed(119, D_WIDTH),
        to_signed(123, D_WIDTH),
        to_signed(126, D_WIDTH),
        to_signed(129, D_WIDTH),
        to_signed(132, D_WIDTH),
        to_signed(136, D_WIDTH),
        to_signed(139, D_WIDTH),
        to_signed(142, D_WIDTH),
        to_signed(145, D_WIDTH),
        to_signed(148, D_WIDTH),
        to_signed(151, D_WIDTH),
        to_signed(154, D_WIDTH),
        to_signed(157, D_WIDTH),
        to_signed(160, D_WIDTH),
        to_signed(163, D_WIDTH),
        to_signed(165, D_WIDTH),
        to_signed(168, D_WIDTH),
        to_signed(171, D_WIDTH),
        to_signed(174, D_WIDTH),
        to_signed(176, D_WIDTH),
        to_signed(179, D_WIDTH),
        to_signed(181, D_WIDTH),
        to_signed(184, D_WIDTH),
        to_signed(186, D_WIDTH),
        to_signed(189, D_WIDTH),
        to_signed(191, D_WIDTH),
        to_signed(193, D_WIDTH),
        to_signed(195, D_WIDTH),
        to_signed(198, D_WIDTH),
        to_signed(200, D_WIDTH),
        to_signed(202, D_WIDTH),
        to_signed(204, D_WIDTH),
        to_signed(206, D_WIDTH),
        to_signed(208, D_WIDTH),
        to_signed(209, D_WIDTH),
        to_signed(211, D_WIDTH),
        to_signed(213, D_WIDTH),
        to_signed(214, D_WIDTH),
        to_signed(216, D_WIDTH),
        to_signed(217, D_WIDTH),
        to_signed(219, D_WIDTH),
        to_signed(220, D_WIDTH),
        to_signed(221, D_WIDTH),
        to_signed(223, D_WIDTH),
        to_signed(224, D_WIDTH),
        to_signed(225, D_WIDTH),
        to_signed(226, D_WIDTH),
        to_signed(227, D_WIDTH),
        to_signed(228, D_WIDTH),
        to_signed(229, D_WIDTH),
        to_signed(229, D_WIDTH),
        to_signed(230, D_WIDTH),
        to_signed(230, D_WIDTH),
        to_signed(231, D_WIDTH),
        to_signed(231, D_WIDTH),
        to_signed(232, D_WIDTH),
        to_signed(232, D_WIDTH),
        to_signed(232, D_WIDTH),
        to_signed(232, D_WIDTH),
        to_signed(232, D_WIDTH),
        to_signed(232, D_WIDTH),
        to_signed(232, D_WIDTH),
        to_signed(232, D_WIDTH),
        to_signed(232, D_WIDTH),
        to_signed(231, D_WIDTH),
        to_signed(231, D_WIDTH),
        to_signed(230, D_WIDTH),
        to_signed(230, D_WIDTH),
        to_signed(229, D_WIDTH),
        to_signed(228, D_WIDTH),
        to_signed(227, D_WIDTH),
        to_signed(226, D_WIDTH),
        to_signed(225, D_WIDTH),
        to_signed(224, D_WIDTH),
        to_signed(223, D_WIDTH),
        to_signed(222, D_WIDTH),
        to_signed(220, D_WIDTH),
        to_signed(219, D_WIDTH),
        to_signed(217, D_WIDTH),
        to_signed(216, D_WIDTH),
        to_signed(214, D_WIDTH),
        to_signed(212, D_WIDTH),
        to_signed(211, D_WIDTH),
        to_signed(209, D_WIDTH),
        to_signed(207, D_WIDTH),
        to_signed(205, D_WIDTH),
        to_signed(202, D_WIDTH),
        to_signed(200, D_WIDTH),
        to_signed(198, D_WIDTH),
        to_signed(195, D_WIDTH),
        to_signed(193, D_WIDTH),
        to_signed(190, D_WIDTH),
        to_signed(188, D_WIDTH),
        to_signed(185, D_WIDTH),
        to_signed(182, D_WIDTH),
        to_signed(179, D_WIDTH),
        to_signed(176, D_WIDTH),
        to_signed(173, D_WIDTH),
        to_signed(170, D_WIDTH),
        to_signed(167, D_WIDTH),
        to_signed(163, D_WIDTH),
        to_signed(160, D_WIDTH),
        to_signed(156, D_WIDTH),
        to_signed(153, D_WIDTH),
        to_signed(149, D_WIDTH),
        to_signed(146, D_WIDTH),
        to_signed(142, D_WIDTH),
        to_signed(138, D_WIDTH),
        to_signed(134, D_WIDTH),
        to_signed(130, D_WIDTH),
        to_signed(126, D_WIDTH),
        to_signed(122, D_WIDTH),
        to_signed(118, D_WIDTH),
        to_signed(114, D_WIDTH),
        to_signed(109, D_WIDTH),
        to_signed(105, D_WIDTH),
        to_signed(101, D_WIDTH),
        to_signed(96, D_WIDTH),
        to_signed(92, D_WIDTH),
        to_signed(87, D_WIDTH),
        to_signed(82, D_WIDTH),
        to_signed(78, D_WIDTH),
        to_signed(73, D_WIDTH),
        to_signed(68, D_WIDTH),
        to_signed(63, D_WIDTH),
        to_signed(58, D_WIDTH),
        to_signed(53, D_WIDTH),
        to_signed(48, D_WIDTH),
        to_signed(43, D_WIDTH),
        to_signed(38, D_WIDTH),
        to_signed(33, D_WIDTH),
        to_signed(27, D_WIDTH),
        to_signed(22, D_WIDTH),
        to_signed(17, D_WIDTH),
        to_signed(11, D_WIDTH),
        to_signed(6, D_WIDTH),
        to_signed(1, D_WIDTH),
        to_signed(-5, D_WIDTH),
        to_signed(-10, D_WIDTH),
        to_signed(-16, D_WIDTH),
        to_signed(-21, D_WIDTH),
        to_signed(-27, D_WIDTH),
        to_signed(-33, D_WIDTH),
        to_signed(-38, D_WIDTH),
        to_signed(-44, D_WIDTH),
        to_signed(-50, D_WIDTH),
        to_signed(-55, D_WIDTH),
        to_signed(-61, D_WIDTH),
        to_signed(-67, D_WIDTH),
        to_signed(-73, D_WIDTH),
        to_signed(-78, D_WIDTH),
        to_signed(-84, D_WIDTH),
        to_signed(-90, D_WIDTH),
        to_signed(-96, D_WIDTH),
        to_signed(-102, D_WIDTH),
        to_signed(-107, D_WIDTH),
        to_signed(-113, D_WIDTH),
        to_signed(-119, D_WIDTH),
        to_signed(-125, D_WIDTH),
        to_signed(-131, D_WIDTH),
        to_signed(-136, D_WIDTH),
        to_signed(-142, D_WIDTH),
        to_signed(-148, D_WIDTH),
        to_signed(-154, D_WIDTH),
        to_signed(-159, D_WIDTH),
        to_signed(-165, D_WIDTH),
        to_signed(-171, D_WIDTH),
        to_signed(-176, D_WIDTH),
        to_signed(-182, D_WIDTH),
        to_signed(-188, D_WIDTH),
        to_signed(-193, D_WIDTH),
        to_signed(-199, D_WIDTH),
        to_signed(-204, D_WIDTH),
        to_signed(-210, D_WIDTH),
        to_signed(-215, D_WIDTH),
        to_signed(-221, D_WIDTH),
        to_signed(-226, D_WIDTH),
        to_signed(-231, D_WIDTH),
        to_signed(-237, D_WIDTH),
        to_signed(-242, D_WIDTH),
        to_signed(-247, D_WIDTH),
        to_signed(-252, D_WIDTH),
        to_signed(-257, D_WIDTH),
        to_signed(-262, D_WIDTH),
        to_signed(-267, D_WIDTH),
        to_signed(-272, D_WIDTH),
        to_signed(-277, D_WIDTH),
        to_signed(-282, D_WIDTH),
        to_signed(-287, D_WIDTH),
        to_signed(-291, D_WIDTH),
        to_signed(-296, D_WIDTH),
        to_signed(-300, D_WIDTH),
        to_signed(-305, D_WIDTH),
        to_signed(-309, D_WIDTH),
        to_signed(-314, D_WIDTH),
        to_signed(-318, D_WIDTH),
        to_signed(-322, D_WIDTH),
        to_signed(-326, D_WIDTH),
        to_signed(-330, D_WIDTH),
        to_signed(-334, D_WIDTH),
        to_signed(-337, D_WIDTH),
        to_signed(-341, D_WIDTH),
        to_signed(-345, D_WIDTH),
        to_signed(-348, D_WIDTH),
        to_signed(-351, D_WIDTH),
        to_signed(-355, D_WIDTH),
        to_signed(-358, D_WIDTH),
        to_signed(-361, D_WIDTH),
        to_signed(-364, D_WIDTH),
        to_signed(-367, D_WIDTH),
        to_signed(-369, D_WIDTH),
        to_signed(-372, D_WIDTH),
        to_signed(-375, D_WIDTH),
        to_signed(-377, D_WIDTH),
        to_signed(-379, D_WIDTH),
        to_signed(-381, D_WIDTH),
        to_signed(-384, D_WIDTH),
        to_signed(-385, D_WIDTH),
        to_signed(-387, D_WIDTH),
        to_signed(-389, D_WIDTH),
        to_signed(-390, D_WIDTH),
        to_signed(-392, D_WIDTH),
        to_signed(-393, D_WIDTH),
        to_signed(-394, D_WIDTH),
        to_signed(-395, D_WIDTH),
        to_signed(-396, D_WIDTH),
        to_signed(-397, D_WIDTH),
        to_signed(-398, D_WIDTH),
        to_signed(-398, D_WIDTH),
        to_signed(-398, D_WIDTH),
        to_signed(-399, D_WIDTH),
        to_signed(-399, D_WIDTH),
        to_signed(-399, D_WIDTH),
        to_signed(-399, D_WIDTH),
        to_signed(-398, D_WIDTH),
        to_signed(-398, D_WIDTH),
        to_signed(-397, D_WIDTH),
        to_signed(-396, D_WIDTH),
        to_signed(-395, D_WIDTH),
        to_signed(-394, D_WIDTH),
        to_signed(-393, D_WIDTH),
        to_signed(-392, D_WIDTH),
        to_signed(-390, D_WIDTH),
        to_signed(-388, D_WIDTH),
        to_signed(-387, D_WIDTH),
        to_signed(-385, D_WIDTH),
        to_signed(-383, D_WIDTH),
        to_signed(-380, D_WIDTH),
        to_signed(-378, D_WIDTH),
        to_signed(-375, D_WIDTH),
        to_signed(-373, D_WIDTH),
        to_signed(-370, D_WIDTH),
        to_signed(-367, D_WIDTH),
        to_signed(-363, D_WIDTH),
        to_signed(-360, D_WIDTH),
        to_signed(-357, D_WIDTH),
        to_signed(-353, D_WIDTH),
        to_signed(-349, D_WIDTH),
        to_signed(-345, D_WIDTH),
        to_signed(-341, D_WIDTH),
        to_signed(-337, D_WIDTH),
        to_signed(-333, D_WIDTH),
        to_signed(-328, D_WIDTH),
        to_signed(-323, D_WIDTH),
        to_signed(-319, D_WIDTH),
        to_signed(-314, D_WIDTH),
        to_signed(-309, D_WIDTH),
        to_signed(-303, D_WIDTH),
        to_signed(-298, D_WIDTH),
        to_signed(-292, D_WIDTH),
        to_signed(-287, D_WIDTH),
        to_signed(-281, D_WIDTH),
        to_signed(-275, D_WIDTH),
        to_signed(-269, D_WIDTH),
        to_signed(-262, D_WIDTH),
        to_signed(-256, D_WIDTH),
        to_signed(-250, D_WIDTH),
        to_signed(-243, D_WIDTH),
        to_signed(-236, D_WIDTH),
        to_signed(-229, D_WIDTH),
        to_signed(-222, D_WIDTH),
        to_signed(-215, D_WIDTH),
        to_signed(-208, D_WIDTH),
        to_signed(-200, D_WIDTH),
        to_signed(-193, D_WIDTH),
        to_signed(-185, D_WIDTH),
        to_signed(-177, D_WIDTH),
        to_signed(-169, D_WIDTH),
        to_signed(-161, D_WIDTH),
        to_signed(-153, D_WIDTH),
        to_signed(-145, D_WIDTH),
        to_signed(-137, D_WIDTH),
        to_signed(-128, D_WIDTH),
        to_signed(-120, D_WIDTH),
        to_signed(-111, D_WIDTH),
        to_signed(-102, D_WIDTH),
        to_signed(-93, D_WIDTH),
        to_signed(-84, D_WIDTH),
        to_signed(-75, D_WIDTH),
        to_signed(-66, D_WIDTH),
        to_signed(-57, D_WIDTH),
        to_signed(-47, D_WIDTH),
        to_signed(-38, D_WIDTH),
        to_signed(-29, D_WIDTH),
        to_signed(-19, D_WIDTH),
        to_signed(-9, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(10, D_WIDTH),
        to_signed(20, D_WIDTH),
        to_signed(30, D_WIDTH),
        to_signed(40, D_WIDTH),
        to_signed(50, D_WIDTH),
        to_signed(60, D_WIDTH),
        to_signed(70, D_WIDTH),
        to_signed(80, D_WIDTH),
        to_signed(90, D_WIDTH),
        to_signed(100, D_WIDTH),
        to_signed(111, D_WIDTH),
        to_signed(121, D_WIDTH),
        to_signed(131, D_WIDTH),
        to_signed(142, D_WIDTH),
        to_signed(152, D_WIDTH),
        to_signed(162, D_WIDTH),
        to_signed(173, D_WIDTH),
        to_signed(183, D_WIDTH),
        to_signed(194, D_WIDTH),
        to_signed(204, D_WIDTH),
        to_signed(214, D_WIDTH),
        to_signed(225, D_WIDTH),
        to_signed(235, D_WIDTH),
        to_signed(246, D_WIDTH),
        to_signed(256, D_WIDTH),
        to_signed(266, D_WIDTH),
        to_signed(277, D_WIDTH),
        to_signed(287, D_WIDTH),
        to_signed(297, D_WIDTH),
        to_signed(307, D_WIDTH),
        to_signed(318, D_WIDTH),
        to_signed(328, D_WIDTH),
        to_signed(338, D_WIDTH),
        to_signed(348, D_WIDTH),
        to_signed(358, D_WIDTH),
        to_signed(368, D_WIDTH),
        to_signed(378, D_WIDTH),
        to_signed(388, D_WIDTH),
        to_signed(397, D_WIDTH),
        to_signed(407, D_WIDTH),
        to_signed(417, D_WIDTH),
        to_signed(426, D_WIDTH),
        to_signed(436, D_WIDTH),
        to_signed(445, D_WIDTH),
        to_signed(454, D_WIDTH),
        to_signed(463, D_WIDTH),
        to_signed(472, D_WIDTH),
        to_signed(481, D_WIDTH),
        to_signed(490, D_WIDTH),
        to_signed(499, D_WIDTH),
        to_signed(507, D_WIDTH),
        to_signed(516, D_WIDTH),
        to_signed(524, D_WIDTH),
        to_signed(532, D_WIDTH),
        to_signed(540, D_WIDTH),
        to_signed(548, D_WIDTH),
        to_signed(556, D_WIDTH),
        to_signed(564, D_WIDTH),
        to_signed(571, D_WIDTH),
        to_signed(579, D_WIDTH),
        to_signed(586, D_WIDTH),
        to_signed(593, D_WIDTH),
        to_signed(600, D_WIDTH),
        to_signed(606, D_WIDTH),
        to_signed(613, D_WIDTH),
        to_signed(619, D_WIDTH),
        to_signed(625, D_WIDTH),
        to_signed(631, D_WIDTH),
        to_signed(637, D_WIDTH),
        to_signed(643, D_WIDTH),
        to_signed(648, D_WIDTH),
        to_signed(654, D_WIDTH),
        to_signed(659, D_WIDTH),
        to_signed(663, D_WIDTH),
        to_signed(668, D_WIDTH),
        to_signed(673, D_WIDTH),
        to_signed(677, D_WIDTH),
        to_signed(681, D_WIDTH),
        to_signed(685, D_WIDTH),
        to_signed(688, D_WIDTH),
        to_signed(691, D_WIDTH),
        to_signed(695, D_WIDTH),
        to_signed(698, D_WIDTH),
        to_signed(700, D_WIDTH),
        to_signed(703, D_WIDTH),
        to_signed(705, D_WIDTH),
        to_signed(707, D_WIDTH),
        to_signed(709, D_WIDTH),
        to_signed(710, D_WIDTH),
        to_signed(711, D_WIDTH),
        to_signed(712, D_WIDTH),
        to_signed(713, D_WIDTH),
        to_signed(714, D_WIDTH),
        to_signed(714, D_WIDTH),
        to_signed(714, D_WIDTH),
        to_signed(714, D_WIDTH),
        to_signed(713, D_WIDTH),
        to_signed(712, D_WIDTH),
        to_signed(711, D_WIDTH),
        to_signed(710, D_WIDTH),
        to_signed(709, D_WIDTH),
        to_signed(707, D_WIDTH),
        to_signed(705, D_WIDTH),
        to_signed(702, D_WIDTH),
        to_signed(700, D_WIDTH),
        to_signed(697, D_WIDTH),
        to_signed(694, D_WIDTH),
        to_signed(690, D_WIDTH),
        to_signed(687, D_WIDTH),
        to_signed(683, D_WIDTH),
        to_signed(679, D_WIDTH),
        to_signed(674, D_WIDTH),
        to_signed(670, D_WIDTH),
        to_signed(665, D_WIDTH),
        to_signed(659, D_WIDTH),
        to_signed(654, D_WIDTH),
        to_signed(648, D_WIDTH),
        to_signed(642, D_WIDTH),
        to_signed(635, D_WIDTH),
        to_signed(629, D_WIDTH),
        to_signed(622, D_WIDTH),
        to_signed(615, D_WIDTH),
        to_signed(607, D_WIDTH),
        to_signed(600, D_WIDTH),
        to_signed(592, D_WIDTH),
        to_signed(584, D_WIDTH),
        to_signed(575, D_WIDTH),
        to_signed(566, D_WIDTH),
        to_signed(557, D_WIDTH),
        to_signed(548, D_WIDTH),
        to_signed(539, D_WIDTH),
        to_signed(529, D_WIDTH),
        to_signed(519, D_WIDTH),
        to_signed(509, D_WIDTH),
        to_signed(498, D_WIDTH),
        to_signed(487, D_WIDTH),
        to_signed(476, D_WIDTH),
        to_signed(465, D_WIDTH),
        to_signed(454, D_WIDTH),
        to_signed(442, D_WIDTH),
        to_signed(430, D_WIDTH),
        to_signed(418, D_WIDTH),
        to_signed(406, D_WIDTH),
        to_signed(393, D_WIDTH),
        to_signed(380, D_WIDTH),
        to_signed(367, D_WIDTH),
        to_signed(354, D_WIDTH),
        to_signed(340, D_WIDTH),
        to_signed(327, D_WIDTH),
        to_signed(313, D_WIDTH),
        to_signed(299, D_WIDTH),
        to_signed(284, D_WIDTH),
        to_signed(270, D_WIDTH),
        to_signed(255, D_WIDTH),
        to_signed(240, D_WIDTH),
        to_signed(225, D_WIDTH),
        to_signed(210, D_WIDTH),
        to_signed(195, D_WIDTH),
        to_signed(179, D_WIDTH),
        to_signed(163, D_WIDTH),
        to_signed(148, D_WIDTH),
        to_signed(132, D_WIDTH),
        to_signed(115, D_WIDTH),
        to_signed(99, D_WIDTH),
        to_signed(83, D_WIDTH),
        to_signed(66, D_WIDTH),
        to_signed(49, D_WIDTH),
        to_signed(32, D_WIDTH),
        to_signed(15, D_WIDTH),
        to_signed(-2, D_WIDTH),
        to_signed(-19, D_WIDTH),
        to_signed(-36, D_WIDTH),
        to_signed(-54, D_WIDTH),
        to_signed(-71, D_WIDTH),
        to_signed(-89, D_WIDTH),
        to_signed(-106, D_WIDTH),
        to_signed(-124, D_WIDTH),
        to_signed(-142, D_WIDTH),
        to_signed(-160, D_WIDTH),
        to_signed(-178, D_WIDTH),
        to_signed(-196, D_WIDTH),
        to_signed(-214, D_WIDTH),
        to_signed(-232, D_WIDTH),
        to_signed(-250, D_WIDTH),
        to_signed(-268, D_WIDTH),
        to_signed(-286, D_WIDTH),
        to_signed(-304, D_WIDTH),
        to_signed(-322, D_WIDTH),
        to_signed(-340, D_WIDTH),
        to_signed(-359, D_WIDTH),
        to_signed(-377, D_WIDTH),
        to_signed(-395, D_WIDTH),
        to_signed(-413, D_WIDTH),
        to_signed(-431, D_WIDTH),
        to_signed(-449, D_WIDTH),
        to_signed(-467, D_WIDTH),
        to_signed(-485, D_WIDTH),
        to_signed(-503, D_WIDTH),
        to_signed(-520, D_WIDTH),
        to_signed(-538, D_WIDTH),
        to_signed(-556, D_WIDTH),
        to_signed(-573, D_WIDTH),
        to_signed(-591, D_WIDTH),
        to_signed(-608, D_WIDTH),
        to_signed(-625, D_WIDTH),
        to_signed(-643, D_WIDTH),
        to_signed(-660, D_WIDTH),
        to_signed(-676, D_WIDTH),
        to_signed(-693, D_WIDTH),
        to_signed(-710, D_WIDTH),
        to_signed(-726, D_WIDTH),
        to_signed(-743, D_WIDTH),
        to_signed(-759, D_WIDTH),
        to_signed(-775, D_WIDTH),
        to_signed(-790, D_WIDTH),
        to_signed(-806, D_WIDTH),
        to_signed(-822, D_WIDTH),
        to_signed(-837, D_WIDTH),
        to_signed(-852, D_WIDTH),
        to_signed(-867, D_WIDTH),
        to_signed(-881, D_WIDTH),
        to_signed(-896, D_WIDTH),
        to_signed(-910, D_WIDTH),
        to_signed(-924, D_WIDTH),
        to_signed(-937, D_WIDTH),
        to_signed(-951, D_WIDTH),
        to_signed(-964, D_WIDTH),
        to_signed(-977, D_WIDTH),
        to_signed(-990, D_WIDTH),
        to_signed(-1002, D_WIDTH),
        to_signed(-1014, D_WIDTH),
        to_signed(-1026, D_WIDTH),
        to_signed(-1037, D_WIDTH),
        to_signed(-1049, D_WIDTH),
        to_signed(-1059, D_WIDTH),
        to_signed(-1070, D_WIDTH),
        to_signed(-1080, D_WIDTH),
        to_signed(-1090, D_WIDTH),
        to_signed(-1100, D_WIDTH),
        to_signed(-1109, D_WIDTH),
        to_signed(-1118, D_WIDTH),
        to_signed(-1127, D_WIDTH),
        to_signed(-1135, D_WIDTH),
        to_signed(-1143, D_WIDTH),
        to_signed(-1151, D_WIDTH),
        to_signed(-1158, D_WIDTH),
        to_signed(-1165, D_WIDTH),
        to_signed(-1171, D_WIDTH),
        to_signed(-1178, D_WIDTH),
        to_signed(-1183, D_WIDTH),
        to_signed(-1189, D_WIDTH),
        to_signed(-1194, D_WIDTH),
        to_signed(-1198, D_WIDTH),
        to_signed(-1202, D_WIDTH),
        to_signed(-1206, D_WIDTH),
        to_signed(-1210, D_WIDTH),
        to_signed(-1213, D_WIDTH),
        to_signed(-1215, D_WIDTH),
        to_signed(-1217, D_WIDTH),
        to_signed(-1219, D_WIDTH),
        to_signed(-1220, D_WIDTH),
        to_signed(-1221, D_WIDTH),
        to_signed(-1222, D_WIDTH),
        to_signed(-1222, D_WIDTH),
        to_signed(-1221, D_WIDTH),
        to_signed(-1221, D_WIDTH),
        to_signed(-1219, D_WIDTH),
        to_signed(-1218, D_WIDTH),
        to_signed(-1215, D_WIDTH),
        to_signed(-1213, D_WIDTH),
        to_signed(-1210, D_WIDTH),
        to_signed(-1206, D_WIDTH),
        to_signed(-1202, D_WIDTH),
        to_signed(-1198, D_WIDTH),
        to_signed(-1193, D_WIDTH),
        to_signed(-1188, D_WIDTH),
        to_signed(-1182, D_WIDTH),
        to_signed(-1176, D_WIDTH),
        to_signed(-1169, D_WIDTH),
        to_signed(-1162, D_WIDTH),
        to_signed(-1155, D_WIDTH),
        to_signed(-1147, D_WIDTH),
        to_signed(-1138, D_WIDTH),
        to_signed(-1129, D_WIDTH),
        to_signed(-1120, D_WIDTH),
        to_signed(-1110, D_WIDTH),
        to_signed(-1100, D_WIDTH),
        to_signed(-1089, D_WIDTH),
        to_signed(-1078, D_WIDTH),
        to_signed(-1067, D_WIDTH),
        to_signed(-1055, D_WIDTH),
        to_signed(-1042, D_WIDTH),
        to_signed(-1029, D_WIDTH),
        to_signed(-1016, D_WIDTH),
        to_signed(-1002, D_WIDTH),
        to_signed(-988, D_WIDTH),
        to_signed(-973, D_WIDTH),
        to_signed(-958, D_WIDTH),
        to_signed(-943, D_WIDTH),
        to_signed(-927, D_WIDTH),
        to_signed(-910, D_WIDTH),
        to_signed(-893, D_WIDTH),
        to_signed(-876, D_WIDTH),
        to_signed(-859, D_WIDTH),
        to_signed(-841, D_WIDTH),
        to_signed(-822, D_WIDTH),
        to_signed(-803, D_WIDTH),
        to_signed(-784, D_WIDTH),
        to_signed(-765, D_WIDTH),
        to_signed(-745, D_WIDTH),
        to_signed(-724, D_WIDTH),
        to_signed(-704, D_WIDTH),
        to_signed(-682, D_WIDTH),
        to_signed(-661, D_WIDTH),
        to_signed(-639, D_WIDTH),
        to_signed(-617, D_WIDTH),
        to_signed(-594, D_WIDTH),
        to_signed(-572, D_WIDTH),
        to_signed(-548, D_WIDTH),
        to_signed(-525, D_WIDTH),
        to_signed(-501, D_WIDTH),
        to_signed(-477, D_WIDTH),
        to_signed(-452, D_WIDTH),
        to_signed(-428, D_WIDTH),
        to_signed(-403, D_WIDTH),
        to_signed(-377, D_WIDTH),
        to_signed(-352, D_WIDTH),
        to_signed(-326, D_WIDTH),
        to_signed(-300, D_WIDTH),
        to_signed(-273, D_WIDTH),
        to_signed(-246, D_WIDTH),
        to_signed(-220, D_WIDTH),
        to_signed(-192, D_WIDTH),
        to_signed(-165, D_WIDTH),
        to_signed(-137, D_WIDTH),
        to_signed(-110, D_WIDTH),
        to_signed(-82, D_WIDTH),
        to_signed(-54, D_WIDTH),
        to_signed(-25, D_WIDTH),
        to_signed(3, D_WIDTH),
        to_signed(32, D_WIDTH),
        to_signed(61, D_WIDTH),
        to_signed(90, D_WIDTH),
        to_signed(119, D_WIDTH),
        to_signed(148, D_WIDTH),
        to_signed(178, D_WIDTH),
        to_signed(207, D_WIDTH),
        to_signed(237, D_WIDTH),
        to_signed(266, D_WIDTH),
        to_signed(296, D_WIDTH),
        to_signed(326, D_WIDTH),
        to_signed(356, D_WIDTH),
        to_signed(385, D_WIDTH),
        to_signed(415, D_WIDTH),
        to_signed(445, D_WIDTH),
        to_signed(475, D_WIDTH),
        to_signed(505, D_WIDTH),
        to_signed(535, D_WIDTH),
        to_signed(565, D_WIDTH),
        to_signed(595, D_WIDTH),
        to_signed(625, D_WIDTH),
        to_signed(655, D_WIDTH),
        to_signed(684, D_WIDTH),
        to_signed(714, D_WIDTH),
        to_signed(744, D_WIDTH),
        to_signed(773, D_WIDTH),
        to_signed(802, D_WIDTH),
        to_signed(832, D_WIDTH),
        to_signed(861, D_WIDTH),
        to_signed(890, D_WIDTH),
        to_signed(919, D_WIDTH),
        to_signed(947, D_WIDTH),
        to_signed(976, D_WIDTH),
        to_signed(1004, D_WIDTH),
        to_signed(1032, D_WIDTH),
        to_signed(1060, D_WIDTH),
        to_signed(1088, D_WIDTH),
        to_signed(1116, D_WIDTH),
        to_signed(1143, D_WIDTH),
        to_signed(1170, D_WIDTH),
        to_signed(1197, D_WIDTH),
        to_signed(1223, D_WIDTH),
        to_signed(1249, D_WIDTH),
        to_signed(1275, D_WIDTH),
        to_signed(1301, D_WIDTH),
        to_signed(1326, D_WIDTH),
        to_signed(1351, D_WIDTH),
        to_signed(1375, D_WIDTH),
        to_signed(1400, D_WIDTH),
        to_signed(1424, D_WIDTH),
        to_signed(1447, D_WIDTH),
        to_signed(1470, D_WIDTH),
        to_signed(1493, D_WIDTH),
        to_signed(1515, D_WIDTH),
        to_signed(1537, D_WIDTH),
        to_signed(1559, D_WIDTH),
        to_signed(1580, D_WIDTH),
        to_signed(1601, D_WIDTH),
        to_signed(1621, D_WIDTH),
        to_signed(1641, D_WIDTH),
        to_signed(1660, D_WIDTH),
        to_signed(1679, D_WIDTH),
        to_signed(1697, D_WIDTH),
        to_signed(1715, D_WIDTH),
        to_signed(1732, D_WIDTH),
        to_signed(1749, D_WIDTH),
        to_signed(1765, D_WIDTH),
        to_signed(1781, D_WIDTH),
        to_signed(1796, D_WIDTH),
        to_signed(1811, D_WIDTH),
        to_signed(1825, D_WIDTH),
        to_signed(1839, D_WIDTH),
        to_signed(1852, D_WIDTH),
        to_signed(1864, D_WIDTH),
        to_signed(1876, D_WIDTH),
        to_signed(1887, D_WIDTH),
        to_signed(1898, D_WIDTH),
        to_signed(1908, D_WIDTH),
        to_signed(1917, D_WIDTH),
        to_signed(1926, D_WIDTH),
        to_signed(1934, D_WIDTH),
        to_signed(1942, D_WIDTH),
        to_signed(1949, D_WIDTH),
        to_signed(1955, D_WIDTH),
        to_signed(1960, D_WIDTH),
        to_signed(1965, D_WIDTH),
        to_signed(1970, D_WIDTH),
        to_signed(1973, D_WIDTH),
        to_signed(1976, D_WIDTH),
        to_signed(1978, D_WIDTH),
        to_signed(1980, D_WIDTH),
        to_signed(1981, D_WIDTH),
        to_signed(1981, D_WIDTH),
        to_signed(1980, D_WIDTH),
        to_signed(1979, D_WIDTH),
        to_signed(1977, D_WIDTH),
        to_signed(1975, D_WIDTH),
        to_signed(1971, D_WIDTH),
        to_signed(1967, D_WIDTH),
        to_signed(1962, D_WIDTH),
        to_signed(1957, D_WIDTH),
        to_signed(1951, D_WIDTH),
        to_signed(1944, D_WIDTH),
        to_signed(1936, D_WIDTH),
        to_signed(1928, D_WIDTH),
        to_signed(1919, D_WIDTH),
        to_signed(1909, D_WIDTH),
        to_signed(1899, D_WIDTH),
        to_signed(1887, D_WIDTH),
        to_signed(1875, D_WIDTH),
        to_signed(1863, D_WIDTH),
        to_signed(1849, D_WIDTH),
        to_signed(1835, D_WIDTH),
        to_signed(1820, D_WIDTH),
        to_signed(1805, D_WIDTH),
        to_signed(1788, D_WIDTH),
        to_signed(1771, D_WIDTH),
        to_signed(1754, D_WIDTH),
        to_signed(1735, D_WIDTH),
        to_signed(1716, D_WIDTH),
        to_signed(1696, D_WIDTH),
        to_signed(1676, D_WIDTH),
        to_signed(1655, D_WIDTH),
        to_signed(1633, D_WIDTH),
        to_signed(1610, D_WIDTH),
        to_signed(1587, D_WIDTH),
        to_signed(1563, D_WIDTH),
        to_signed(1538, D_WIDTH),
        to_signed(1513, D_WIDTH),
        to_signed(1487, D_WIDTH),
        to_signed(1460, D_WIDTH),
        to_signed(1433, D_WIDTH),
        to_signed(1405, D_WIDTH),
        to_signed(1376, D_WIDTH),
        to_signed(1347, D_WIDTH),
        to_signed(1317, D_WIDTH),
        to_signed(1287, D_WIDTH),
        to_signed(1256, D_WIDTH),
        to_signed(1224, D_WIDTH),
        to_signed(1192, D_WIDTH),
        to_signed(1159, D_WIDTH),
        to_signed(1126, D_WIDTH),
        to_signed(1092, D_WIDTH),
        to_signed(1057, D_WIDTH),
        to_signed(1022, D_WIDTH),
        to_signed(986, D_WIDTH),
        to_signed(950, D_WIDTH),
        to_signed(913, D_WIDTH),
        to_signed(876, D_WIDTH),
        to_signed(838, D_WIDTH),
        to_signed(800, D_WIDTH),
        to_signed(761, D_WIDTH),
        to_signed(722, D_WIDTH),
        to_signed(682, D_WIDTH),
        to_signed(642, D_WIDTH),
        to_signed(602, D_WIDTH),
        to_signed(561, D_WIDTH),
        to_signed(519, D_WIDTH),
        to_signed(478, D_WIDTH),
        to_signed(435, D_WIDTH),
        to_signed(393, D_WIDTH),
        to_signed(350, D_WIDTH),
        to_signed(307, D_WIDTH),
        to_signed(263, D_WIDTH),
        to_signed(219, D_WIDTH),
        to_signed(175, D_WIDTH),
        to_signed(131, D_WIDTH),
        to_signed(86, D_WIDTH),
        to_signed(41, D_WIDTH),
        to_signed(-4, D_WIDTH),
        to_signed(-50, D_WIDTH),
        to_signed(-96, D_WIDTH),
        to_signed(-142, D_WIDTH),
        to_signed(-188, D_WIDTH),
        to_signed(-234, D_WIDTH),
        to_signed(-280, D_WIDTH),
        to_signed(-327, D_WIDTH),
        to_signed(-374, D_WIDTH),
        to_signed(-421, D_WIDTH),
        to_signed(-468, D_WIDTH),
        to_signed(-515, D_WIDTH),
        to_signed(-562, D_WIDTH),
        to_signed(-609, D_WIDTH),
        to_signed(-656, D_WIDTH),
        to_signed(-703, D_WIDTH),
        to_signed(-750, D_WIDTH),
        to_signed(-797, D_WIDTH),
        to_signed(-845, D_WIDTH),
        to_signed(-892, D_WIDTH),
        to_signed(-939, D_WIDTH),
        to_signed(-986, D_WIDTH),
        to_signed(-1032, D_WIDTH),
        to_signed(-1079, D_WIDTH),
        to_signed(-1126, D_WIDTH),
        to_signed(-1172, D_WIDTH),
        to_signed(-1218, D_WIDTH),
        to_signed(-1264, D_WIDTH),
        to_signed(-1310, D_WIDTH),
        to_signed(-1356, D_WIDTH),
        to_signed(-1401, D_WIDTH),
        to_signed(-1446, D_WIDTH),
        to_signed(-1491, D_WIDTH),
        to_signed(-1536, D_WIDTH),
        to_signed(-1580, D_WIDTH),
        to_signed(-1624, D_WIDTH),
        to_signed(-1667, D_WIDTH),
        to_signed(-1710, D_WIDTH),
        to_signed(-1753, D_WIDTH),
        to_signed(-1796, D_WIDTH),
        to_signed(-1838, D_WIDTH),
        to_signed(-1879, D_WIDTH),
        to_signed(-1921, D_WIDTH),
        to_signed(-1961, D_WIDTH),
        to_signed(-2001, D_WIDTH),
        to_signed(-2041, D_WIDTH),
        to_signed(-2080, D_WIDTH),
        to_signed(-2119, D_WIDTH),
        to_signed(-2157, D_WIDTH),
        to_signed(-2195, D_WIDTH),
        to_signed(-2232, D_WIDTH),
        to_signed(-2268, D_WIDTH),
        to_signed(-2304, D_WIDTH),
        to_signed(-2339, D_WIDTH),
        to_signed(-2374, D_WIDTH),
        to_signed(-2408, D_WIDTH),
        to_signed(-2441, D_WIDTH),
        to_signed(-2473, D_WIDTH),
        to_signed(-2505, D_WIDTH),
        to_signed(-2536, D_WIDTH),
        to_signed(-2567, D_WIDTH),
        to_signed(-2596, D_WIDTH),
        to_signed(-2625, D_WIDTH),
        to_signed(-2653, D_WIDTH),
        to_signed(-2681, D_WIDTH),
        to_signed(-2707, D_WIDTH),
        to_signed(-2733, D_WIDTH),
        to_signed(-2758, D_WIDTH),
        to_signed(-2782, D_WIDTH),
        to_signed(-2805, D_WIDTH),
        to_signed(-2828, D_WIDTH),
        to_signed(-2849, D_WIDTH),
        to_signed(-2870, D_WIDTH),
        to_signed(-2889, D_WIDTH),
        to_signed(-2908, D_WIDTH),
        to_signed(-2926, D_WIDTH),
        to_signed(-2943, D_WIDTH),
        to_signed(-2959, D_WIDTH),
        to_signed(-2974, D_WIDTH),
        to_signed(-2988, D_WIDTH),
        to_signed(-3001, D_WIDTH),
        to_signed(-3013, D_WIDTH),
        to_signed(-3024, D_WIDTH),
        to_signed(-3034, D_WIDTH),
        to_signed(-3044, D_WIDTH),
        to_signed(-3052, D_WIDTH),
        to_signed(-3059, D_WIDTH),
        to_signed(-3065, D_WIDTH),
        to_signed(-3070, D_WIDTH),
        to_signed(-3074, D_WIDTH),
        to_signed(-3077, D_WIDTH),
        to_signed(-3078, D_WIDTH),
        to_signed(-3079, D_WIDTH),
        to_signed(-3079, D_WIDTH),
        to_signed(-3078, D_WIDTH),
        to_signed(-3075, D_WIDTH),
        to_signed(-3072, D_WIDTH),
        to_signed(-3067, D_WIDTH),
        to_signed(-3061, D_WIDTH),
        to_signed(-3054, D_WIDTH),
        to_signed(-3046, D_WIDTH),
        to_signed(-3037, D_WIDTH),
        to_signed(-3027, D_WIDTH),
        to_signed(-3016, D_WIDTH),
        to_signed(-3004, D_WIDTH),
        to_signed(-2990, D_WIDTH),
        to_signed(-2976, D_WIDTH),
        to_signed(-2960, D_WIDTH),
        to_signed(-2943, D_WIDTH),
        to_signed(-2925, D_WIDTH),
        to_signed(-2906, D_WIDTH),
        to_signed(-2886, D_WIDTH),
        to_signed(-2865, D_WIDTH),
        to_signed(-2842, D_WIDTH),
        to_signed(-2819, D_WIDTH),
        to_signed(-2794, D_WIDTH),
        to_signed(-2769, D_WIDTH),
        to_signed(-2742, D_WIDTH),
        to_signed(-2714, D_WIDTH),
        to_signed(-2685, D_WIDTH),
        to_signed(-2655, D_WIDTH),
        to_signed(-2624, D_WIDTH),
        to_signed(-2592, D_WIDTH),
        to_signed(-2559, D_WIDTH),
        to_signed(-2525, D_WIDTH),
        to_signed(-2489, D_WIDTH),
        to_signed(-2453, D_WIDTH),
        to_signed(-2416, D_WIDTH),
        to_signed(-2377, D_WIDTH),
        to_signed(-2338, D_WIDTH),
        to_signed(-2297, D_WIDTH),
        to_signed(-2256, D_WIDTH),
        to_signed(-2213, D_WIDTH),
        to_signed(-2170, D_WIDTH),
        to_signed(-2125, D_WIDTH),
        to_signed(-2080, D_WIDTH),
        to_signed(-2034, D_WIDTH),
        to_signed(-1986, D_WIDTH),
        to_signed(-1938, D_WIDTH),
        to_signed(-1889, D_WIDTH),
        to_signed(-1839, D_WIDTH),
        to_signed(-1788, D_WIDTH),
        to_signed(-1736, D_WIDTH),
        to_signed(-1684, D_WIDTH),
        to_signed(-1630, D_WIDTH),
        to_signed(-1576, D_WIDTH),
        to_signed(-1521, D_WIDTH),
        to_signed(-1465, D_WIDTH),
        to_signed(-1408, D_WIDTH),
        to_signed(-1351, D_WIDTH),
        to_signed(-1293, D_WIDTH),
        to_signed(-1234, D_WIDTH),
        to_signed(-1174, D_WIDTH),
        to_signed(-1113, D_WIDTH),
        to_signed(-1052, D_WIDTH),
        to_signed(-991, D_WIDTH),
        to_signed(-928, D_WIDTH),
        to_signed(-865, D_WIDTH),
        to_signed(-801, D_WIDTH),
        to_signed(-737, D_WIDTH),
        to_signed(-672, D_WIDTH),
        to_signed(-607, D_WIDTH),
        to_signed(-541, D_WIDTH),
        to_signed(-475, D_WIDTH),
        to_signed(-408, D_WIDTH),
        to_signed(-340, D_WIDTH),
        to_signed(-272, D_WIDTH),
        to_signed(-204, D_WIDTH),
        to_signed(-136, D_WIDTH),
        to_signed(-66, D_WIDTH),
        to_signed(3, D_WIDTH),
        to_signed(73, D_WIDTH),
        to_signed(143, D_WIDTH),
        to_signed(213, D_WIDTH),
        to_signed(284, D_WIDTH),
        to_signed(355, D_WIDTH),
        to_signed(426, D_WIDTH),
        to_signed(497, D_WIDTH),
        to_signed(569, D_WIDTH),
        to_signed(640, D_WIDTH),
        to_signed(712, D_WIDTH),
        to_signed(784, D_WIDTH),
        to_signed(856, D_WIDTH),
        to_signed(928, D_WIDTH),
        to_signed(1000, D_WIDTH),
        to_signed(1072, D_WIDTH),
        to_signed(1144, D_WIDTH),
        to_signed(1216, D_WIDTH),
        to_signed(1288, D_WIDTH),
        to_signed(1360, D_WIDTH),
        to_signed(1431, D_WIDTH),
        to_signed(1503, D_WIDTH),
        to_signed(1574, D_WIDTH),
        to_signed(1646, D_WIDTH),
        to_signed(1717, D_WIDTH),
        to_signed(1787, D_WIDTH),
        to_signed(1858, D_WIDTH),
        to_signed(1928, D_WIDTH),
        to_signed(1998, D_WIDTH),
        to_signed(2067, D_WIDTH),
        to_signed(2136, D_WIDTH),
        to_signed(2205, D_WIDTH),
        to_signed(2273, D_WIDTH),
        to_signed(2341, D_WIDTH),
        to_signed(2408, D_WIDTH),
        to_signed(2475, D_WIDTH),
        to_signed(2541, D_WIDTH),
        to_signed(2607, D_WIDTH),
        to_signed(2672, D_WIDTH),
        to_signed(2736, D_WIDTH),
        to_signed(2800, D_WIDTH),
        to_signed(2863, D_WIDTH),
        to_signed(2926, D_WIDTH),
        to_signed(2987, D_WIDTH),
        to_signed(3048, D_WIDTH),
        to_signed(3109, D_WIDTH),
        to_signed(3168, D_WIDTH),
        to_signed(3227, D_WIDTH),
        to_signed(3285, D_WIDTH),
        to_signed(3342, D_WIDTH),
        to_signed(3398, D_WIDTH),
        to_signed(3453, D_WIDTH),
        to_signed(3507, D_WIDTH),
        to_signed(3560, D_WIDTH),
        to_signed(3613, D_WIDTH),
        to_signed(3664, D_WIDTH),
        to_signed(3714, D_WIDTH),
        to_signed(3763, D_WIDTH),
        to_signed(3812, D_WIDTH),
        to_signed(3859, D_WIDTH),
        to_signed(3905, D_WIDTH),
        to_signed(3949, D_WIDTH),
        to_signed(3993, D_WIDTH),
        to_signed(4035, D_WIDTH),
        to_signed(4077, D_WIDTH),
        to_signed(4117, D_WIDTH),
        to_signed(4156, D_WIDTH),
        to_signed(4193, D_WIDTH),
        to_signed(4229, D_WIDTH),
        to_signed(4264, D_WIDTH),
        to_signed(4298, D_WIDTH),
        to_signed(4330, D_WIDTH),
        to_signed(4361, D_WIDTH),
        to_signed(4391, D_WIDTH),
        to_signed(4419, D_WIDTH),
        to_signed(4446, D_WIDTH),
        to_signed(4472, D_WIDTH),
        to_signed(4496, D_WIDTH),
        to_signed(4518, D_WIDTH),
        to_signed(4539, D_WIDTH),
        to_signed(4559, D_WIDTH),
        to_signed(4577, D_WIDTH),
        to_signed(4593, D_WIDTH),
        to_signed(4609, D_WIDTH),
        to_signed(4622, D_WIDTH),
        to_signed(4634, D_WIDTH),
        to_signed(4645, D_WIDTH),
        to_signed(4653, D_WIDTH),
        to_signed(4661, D_WIDTH),
        to_signed(4667, D_WIDTH),
        to_signed(4671, D_WIDTH),
        to_signed(4673, D_WIDTH),
        to_signed(4674, D_WIDTH),
        to_signed(4673, D_WIDTH),
        to_signed(4671, D_WIDTH),
        to_signed(4667, D_WIDTH),
        to_signed(4662, D_WIDTH),
        to_signed(4654, D_WIDTH),
        to_signed(4645, D_WIDTH),
        to_signed(4635, D_WIDTH),
        to_signed(4623, D_WIDTH),
        to_signed(4609, D_WIDTH),
        to_signed(4593, D_WIDTH),
        to_signed(4576, D_WIDTH),
        to_signed(4557, D_WIDTH),
        to_signed(4536, D_WIDTH),
        to_signed(4514, D_WIDTH),
        to_signed(4490, D_WIDTH),
        to_signed(4464, D_WIDTH),
        to_signed(4437, D_WIDTH),
        to_signed(4408, D_WIDTH),
        to_signed(4377, D_WIDTH),
        to_signed(4345, D_WIDTH),
        to_signed(4311, D_WIDTH),
        to_signed(4275, D_WIDTH),
        to_signed(4238, D_WIDTH),
        to_signed(4199, D_WIDTH),
        to_signed(4158, D_WIDTH),
        to_signed(4116, D_WIDTH),
        to_signed(4072, D_WIDTH),
        to_signed(4027, D_WIDTH),
        to_signed(3980, D_WIDTH),
        to_signed(3931, D_WIDTH),
        to_signed(3880, D_WIDTH),
        to_signed(3828, D_WIDTH),
        to_signed(3775, D_WIDTH),
        to_signed(3720, D_WIDTH),
        to_signed(3663, D_WIDTH),
        to_signed(3605, D_WIDTH),
        to_signed(3545, D_WIDTH),
        to_signed(3484, D_WIDTH),
        to_signed(3421, D_WIDTH),
        to_signed(3356, D_WIDTH),
        to_signed(3291, D_WIDTH),
        to_signed(3223, D_WIDTH),
        to_signed(3155, D_WIDTH),
        to_signed(3085, D_WIDTH),
        to_signed(3013, D_WIDTH),
        to_signed(2940, D_WIDTH),
        to_signed(2866, D_WIDTH),
        to_signed(2790, D_WIDTH),
        to_signed(2713, D_WIDTH),
        to_signed(2635, D_WIDTH),
        to_signed(2555, D_WIDTH),
        to_signed(2474, D_WIDTH),
        to_signed(2392, D_WIDTH),
        to_signed(2308, D_WIDTH),
        to_signed(2224, D_WIDTH),
        to_signed(2138, D_WIDTH),
        to_signed(2051, D_WIDTH),
        to_signed(1963, D_WIDTH),
        to_signed(1874, D_WIDTH),
        to_signed(1783, D_WIDTH),
        to_signed(1692, D_WIDTH),
        to_signed(1600, D_WIDTH),
        to_signed(1506, D_WIDTH),
        to_signed(1412, D_WIDTH),
        to_signed(1317, D_WIDTH),
        to_signed(1220, D_WIDTH),
        to_signed(1123, D_WIDTH),
        to_signed(1025, D_WIDTH),
        to_signed(926, D_WIDTH),
        to_signed(827, D_WIDTH),
        to_signed(726, D_WIDTH),
        to_signed(625, D_WIDTH),
        to_signed(523, D_WIDTH),
        to_signed(420, D_WIDTH),
        to_signed(317, D_WIDTH),
        to_signed(213, D_WIDTH),
        to_signed(109, D_WIDTH),
        to_signed(4, D_WIDTH),
        to_signed(-102, D_WIDTH),
        to_signed(-208, D_WIDTH),
        to_signed(-314, D_WIDTH),
        to_signed(-421, D_WIDTH),
        to_signed(-528, D_WIDTH),
        to_signed(-636, D_WIDTH),
        to_signed(-743, D_WIDTH),
        to_signed(-852, D_WIDTH),
        to_signed(-960, D_WIDTH),
        to_signed(-1069, D_WIDTH),
        to_signed(-1177, D_WIDTH),
        to_signed(-1286, D_WIDTH),
        to_signed(-1395, D_WIDTH),
        to_signed(-1504, D_WIDTH),
        to_signed(-1613, D_WIDTH),
        to_signed(-1722, D_WIDTH),
        to_signed(-1831, D_WIDTH),
        to_signed(-1940, D_WIDTH),
        to_signed(-2048, D_WIDTH),
        to_signed(-2157, D_WIDTH),
        to_signed(-2265, D_WIDTH),
        to_signed(-2373, D_WIDTH),
        to_signed(-2481, D_WIDTH),
        to_signed(-2588, D_WIDTH),
        to_signed(-2696, D_WIDTH),
        to_signed(-2802, D_WIDTH),
        to_signed(-2908, D_WIDTH),
        to_signed(-3014, D_WIDTH),
        to_signed(-3119, D_WIDTH),
        to_signed(-3224, D_WIDTH),
        to_signed(-3328, D_WIDTH),
        to_signed(-3431, D_WIDTH),
        to_signed(-3534, D_WIDTH),
        to_signed(-3636, D_WIDTH),
        to_signed(-3737, D_WIDTH),
        to_signed(-3838, D_WIDTH),
        to_signed(-3937, D_WIDTH),
        to_signed(-4036, D_WIDTH),
        to_signed(-4134, D_WIDTH),
        to_signed(-4230, D_WIDTH),
        to_signed(-4326, D_WIDTH),
        to_signed(-4421, D_WIDTH),
        to_signed(-4515, D_WIDTH),
        to_signed(-4608, D_WIDTH),
        to_signed(-4699, D_WIDTH),
        to_signed(-4789, D_WIDTH),
        to_signed(-4879, D_WIDTH),
        to_signed(-4966, D_WIDTH),
        to_signed(-5053, D_WIDTH),
        to_signed(-5138, D_WIDTH),
        to_signed(-5222, D_WIDTH),
        to_signed(-5305, D_WIDTH),
        to_signed(-5386, D_WIDTH),
        to_signed(-5465, D_WIDTH),
        to_signed(-5543, D_WIDTH),
        to_signed(-5620, D_WIDTH),
        to_signed(-5695, D_WIDTH),
        to_signed(-5768, D_WIDTH),
        to_signed(-5840, D_WIDTH),
        to_signed(-5910, D_WIDTH),
        to_signed(-5979, D_WIDTH),
        to_signed(-6045, D_WIDTH),
        to_signed(-6110, D_WIDTH),
        to_signed(-6173, D_WIDTH),
        to_signed(-6235, D_WIDTH),
        to_signed(-6294, D_WIDTH),
        to_signed(-6351, D_WIDTH),
        to_signed(-6407, D_WIDTH),
        to_signed(-6461, D_WIDTH),
        to_signed(-6512, D_WIDTH),
        to_signed(-6562, D_WIDTH),
        to_signed(-6610, D_WIDTH),
        to_signed(-6655, D_WIDTH),
        to_signed(-6699, D_WIDTH),
        to_signed(-6740, D_WIDTH),
        to_signed(-6780, D_WIDTH),
        to_signed(-6817, D_WIDTH),
        to_signed(-6852, D_WIDTH),
        to_signed(-6884, D_WIDTH),
        to_signed(-6915, D_WIDTH),
        to_signed(-6943, D_WIDTH),
        to_signed(-6969, D_WIDTH),
        to_signed(-6993, D_WIDTH),
        to_signed(-7014, D_WIDTH),
        to_signed(-7033, D_WIDTH),
        to_signed(-7050, D_WIDTH),
        to_signed(-7064, D_WIDTH),
        to_signed(-7076, D_WIDTH),
        to_signed(-7086, D_WIDTH),
        to_signed(-7093, D_WIDTH),
        to_signed(-7098, D_WIDTH),
        to_signed(-7100, D_WIDTH),
        to_signed(-7100, D_WIDTH),
        to_signed(-7098, D_WIDTH),
        to_signed(-7092, D_WIDTH),
        to_signed(-7085, D_WIDTH),
        to_signed(-7075, D_WIDTH),
        to_signed(-7062, D_WIDTH),
        to_signed(-7047, D_WIDTH),
        to_signed(-7030, D_WIDTH),
        to_signed(-7010, D_WIDTH),
        to_signed(-6987, D_WIDTH),
        to_signed(-6962, D_WIDTH),
        to_signed(-6934, D_WIDTH),
        to_signed(-6904, D_WIDTH),
        to_signed(-6871, D_WIDTH),
        to_signed(-6835, D_WIDTH),
        to_signed(-6797, D_WIDTH),
        to_signed(-6757, D_WIDTH),
        to_signed(-6714, D_WIDTH),
        to_signed(-6668, D_WIDTH),
        to_signed(-6620, D_WIDTH),
        to_signed(-6569, D_WIDTH),
        to_signed(-6516, D_WIDTH),
        to_signed(-6460, D_WIDTH),
        to_signed(-6402, D_WIDTH),
        to_signed(-6341, D_WIDTH),
        to_signed(-6278, D_WIDTH),
        to_signed(-6212, D_WIDTH),
        to_signed(-6144, D_WIDTH),
        to_signed(-6073, D_WIDTH),
        to_signed(-6000, D_WIDTH),
        to_signed(-5924, D_WIDTH),
        to_signed(-5846, D_WIDTH),
        to_signed(-5765, D_WIDTH),
        to_signed(-5682, D_WIDTH),
        to_signed(-5597, D_WIDTH),
        to_signed(-5509, D_WIDTH),
        to_signed(-5419, D_WIDTH),
        to_signed(-5326, D_WIDTH),
        to_signed(-5231, D_WIDTH),
        to_signed(-5134, D_WIDTH),
        to_signed(-5035, D_WIDTH),
        to_signed(-4933, D_WIDTH),
        to_signed(-4829, D_WIDTH),
        to_signed(-4723, D_WIDTH),
        to_signed(-4615, D_WIDTH),
        to_signed(-4504, D_WIDTH),
        to_signed(-4391, D_WIDTH),
        to_signed(-4277, D_WIDTH),
        to_signed(-4160, D_WIDTH),
        to_signed(-4041, D_WIDTH),
        to_signed(-3920, D_WIDTH),
        to_signed(-3797, D_WIDTH),
        to_signed(-3672, D_WIDTH),
        to_signed(-3545, D_WIDTH),
        to_signed(-3417, D_WIDTH),
        to_signed(-3286, D_WIDTH),
        to_signed(-3154, D_WIDTH),
        to_signed(-3020, D_WIDTH),
        to_signed(-2884, D_WIDTH),
        to_signed(-2746, D_WIDTH),
        to_signed(-2607, D_WIDTH),
        to_signed(-2466, D_WIDTH),
        to_signed(-2323, D_WIDTH),
        to_signed(-2179, D_WIDTH),
        to_signed(-2033, D_WIDTH),
        to_signed(-1886, D_WIDTH),
        to_signed(-1738, D_WIDTH),
        to_signed(-1588, D_WIDTH),
        to_signed(-1437, D_WIDTH),
        to_signed(-1284, D_WIDTH),
        to_signed(-1130, D_WIDTH),
        to_signed(-975, D_WIDTH),
        to_signed(-819, D_WIDTH),
        to_signed(-662, D_WIDTH),
        to_signed(-503, D_WIDTH),
        to_signed(-344, D_WIDTH),
        to_signed(-183, D_WIDTH),
        to_signed(-22, D_WIDTH),
        to_signed(140, D_WIDTH),
        to_signed(303, D_WIDTH),
        to_signed(467, D_WIDTH),
        to_signed(631, D_WIDTH),
        to_signed(796, D_WIDTH),
        to_signed(962, D_WIDTH),
        to_signed(1128, D_WIDTH),
        to_signed(1295, D_WIDTH),
        to_signed(1463, D_WIDTH),
        to_signed(1630, D_WIDTH),
        to_signed(1798, D_WIDTH),
        to_signed(1966, D_WIDTH),
        to_signed(2135, D_WIDTH),
        to_signed(2304, D_WIDTH),
        to_signed(2472, D_WIDTH),
        to_signed(2641, D_WIDTH),
        to_signed(2810, D_WIDTH),
        to_signed(2979, D_WIDTH),
        to_signed(3147, D_WIDTH),
        to_signed(3316, D_WIDTH),
        to_signed(3484, D_WIDTH),
        to_signed(3652, D_WIDTH),
        to_signed(3820, D_WIDTH),
        to_signed(3987, D_WIDTH),
        to_signed(4154, D_WIDTH),
        to_signed(4320, D_WIDTH),
        to_signed(4486, D_WIDTH),
        to_signed(4651, D_WIDTH),
        to_signed(4815, D_WIDTH),
        to_signed(4978, D_WIDTH),
        to_signed(5141, D_WIDTH),
        to_signed(5303, D_WIDTH),
        to_signed(5464, D_WIDTH),
        to_signed(5624, D_WIDTH),
        to_signed(5782, D_WIDTH),
        to_signed(5940, D_WIDTH),
        to_signed(6096, D_WIDTH),
        to_signed(6252, D_WIDTH),
        to_signed(6406, D_WIDTH),
        to_signed(6558, D_WIDTH),
        to_signed(6709, D_WIDTH),
        to_signed(6859, D_WIDTH),
        to_signed(7007, D_WIDTH),
        to_signed(7154, D_WIDTH),
        to_signed(7298, D_WIDTH),
        to_signed(7441, D_WIDTH),
        to_signed(7583, D_WIDTH),
        to_signed(7722, D_WIDTH),
        to_signed(7860, D_WIDTH),
        to_signed(7996, D_WIDTH),
        to_signed(8129, D_WIDTH),
        to_signed(8261, D_WIDTH),
        to_signed(8390, D_WIDTH),
        to_signed(8517, D_WIDTH),
        to_signed(8643, D_WIDTH),
        to_signed(8765, D_WIDTH),
        to_signed(8886, D_WIDTH),
        to_signed(9004, D_WIDTH),
        to_signed(9119, D_WIDTH),
        to_signed(9232, D_WIDTH),
        to_signed(9343, D_WIDTH),
        to_signed(9451, D_WIDTH),
        to_signed(9556, D_WIDTH),
        to_signed(9658, D_WIDTH),
        to_signed(9758, D_WIDTH),
        to_signed(9855, D_WIDTH),
        to_signed(9949, D_WIDTH),
        to_signed(10040, D_WIDTH),
        to_signed(10129, D_WIDTH),
        to_signed(10214, D_WIDTH),
        to_signed(10296, D_WIDTH),
        to_signed(10375, D_WIDTH),
        to_signed(10451, D_WIDTH),
        to_signed(10524, D_WIDTH),
        to_signed(10593, D_WIDTH),
        to_signed(10660, D_WIDTH),
        to_signed(10723, D_WIDTH),
        to_signed(10782, D_WIDTH),
        to_signed(10838, D_WIDTH),
        to_signed(10891, D_WIDTH),
        to_signed(10940, D_WIDTH),
        to_signed(10986, D_WIDTH),
        to_signed(11029, D_WIDTH),
        to_signed(11067, D_WIDTH),
        to_signed(11102, D_WIDTH),
        to_signed(11134, D_WIDTH),
        to_signed(11162, D_WIDTH),
        to_signed(11186, D_WIDTH),
        to_signed(11206, D_WIDTH),
        to_signed(11223, D_WIDTH),
        to_signed(11235, D_WIDTH),
        to_signed(11244, D_WIDTH),
        to_signed(11249, D_WIDTH),
        to_signed(11251, D_WIDTH),
        to_signed(11248, D_WIDTH),
        to_signed(11242, D_WIDTH),
        to_signed(11231, D_WIDTH),
        to_signed(11217, D_WIDTH),
        to_signed(11198, D_WIDTH),
        to_signed(11176, D_WIDTH),
        to_signed(11149, D_WIDTH),
        to_signed(11119, D_WIDTH),
        to_signed(11084, D_WIDTH),
        to_signed(11046, D_WIDTH),
        to_signed(11003, D_WIDTH),
        to_signed(10957, D_WIDTH),
        to_signed(10906, D_WIDTH),
        to_signed(10851, D_WIDTH),
        to_signed(10792, D_WIDTH),
        to_signed(10729, D_WIDTH),
        to_signed(10662, D_WIDTH),
        to_signed(10591, D_WIDTH),
        to_signed(10515, D_WIDTH),
        to_signed(10436, D_WIDTH),
        to_signed(10353, D_WIDTH),
        to_signed(10265, D_WIDTH),
        to_signed(10173, D_WIDTH),
        to_signed(10077, D_WIDTH),
        to_signed(9977, D_WIDTH),
        to_signed(9873, D_WIDTH),
        to_signed(9765, D_WIDTH),
        to_signed(9653, D_WIDTH),
        to_signed(9537, D_WIDTH),
        to_signed(9417, D_WIDTH),
        to_signed(9293, D_WIDTH),
        to_signed(9164, D_WIDTH),
        to_signed(9032, D_WIDTH),
        to_signed(8896, D_WIDTH),
        to_signed(8756, D_WIDTH),
        to_signed(8612, D_WIDTH),
        to_signed(8464, D_WIDTH),
        to_signed(8312, D_WIDTH),
        to_signed(8157, D_WIDTH),
        to_signed(7997, D_WIDTH),
        to_signed(7834, D_WIDTH),
        to_signed(7667, D_WIDTH),
        to_signed(7497, D_WIDTH),
        to_signed(7322, D_WIDTH),
        to_signed(7144, D_WIDTH),
        to_signed(6963, D_WIDTH),
        to_signed(6777, D_WIDTH),
        to_signed(6589, D_WIDTH),
        to_signed(6396, D_WIDTH),
        to_signed(6201, D_WIDTH),
        to_signed(6002, D_WIDTH),
        to_signed(5799, D_WIDTH),
        to_signed(5593, D_WIDTH),
        to_signed(5384, D_WIDTH),
        to_signed(5172, D_WIDTH),
        to_signed(4956, D_WIDTH),
        to_signed(4738, D_WIDTH),
        to_signed(4516, D_WIDTH),
        to_signed(4291, D_WIDTH),
        to_signed(4064, D_WIDTH),
        to_signed(3833, D_WIDTH),
        to_signed(3600, D_WIDTH),
        to_signed(3363, D_WIDTH),
        to_signed(3124, D_WIDTH),
        to_signed(2883, D_WIDTH),
        to_signed(2638, D_WIDTH),
        to_signed(2392, D_WIDTH),
        to_signed(2142, D_WIDTH),
        to_signed(1891, D_WIDTH),
        to_signed(1637, D_WIDTH),
        to_signed(1380, D_WIDTH),
        to_signed(1122, D_WIDTH),
        to_signed(861, D_WIDTH),
        to_signed(598, D_WIDTH),
        to_signed(334, D_WIDTH),
        to_signed(67, D_WIDTH),
        to_signed(-201, D_WIDTH),
        to_signed(-472, D_WIDTH),
        to_signed(-744, D_WIDTH),
        to_signed(-1017, D_WIDTH),
        to_signed(-1292, D_WIDTH),
        to_signed(-1569, D_WIDTH),
        to_signed(-1847, D_WIDTH),
        to_signed(-2126, D_WIDTH),
        to_signed(-2406, D_WIDTH),
        to_signed(-2688, D_WIDTH),
        to_signed(-2970, D_WIDTH),
        to_signed(-3254, D_WIDTH),
        to_signed(-3538, D_WIDTH),
        to_signed(-3823, D_WIDTH),
        to_signed(-4109, D_WIDTH),
        to_signed(-4395, D_WIDTH),
        to_signed(-4682, D_WIDTH),
        to_signed(-4969, D_WIDTH),
        to_signed(-5257, D_WIDTH),
        to_signed(-5545, D_WIDTH),
        to_signed(-5833, D_WIDTH),
        to_signed(-6121, D_WIDTH),
        to_signed(-6409, D_WIDTH),
        to_signed(-6696, D_WIDTH),
        to_signed(-6984, D_WIDTH),
        to_signed(-7271, D_WIDTH),
        to_signed(-7558, D_WIDTH),
        to_signed(-7844, D_WIDTH),
        to_signed(-8129, D_WIDTH),
        to_signed(-8414, D_WIDTH),
        to_signed(-8698, D_WIDTH),
        to_signed(-8981, D_WIDTH),
        to_signed(-9263, D_WIDTH),
        to_signed(-9544, D_WIDTH),
        to_signed(-9824, D_WIDTH),
        to_signed(-10102, D_WIDTH),
        to_signed(-10379, D_WIDTH),
        to_signed(-10654, D_WIDTH),
        to_signed(-10928, D_WIDTH),
        to_signed(-11200, D_WIDTH),
        to_signed(-11470, D_WIDTH),
        to_signed(-11738, D_WIDTH),
        to_signed(-12004, D_WIDTH),
        to_signed(-12268, D_WIDTH),
        to_signed(-12530, D_WIDTH),
        to_signed(-12789, D_WIDTH),
        to_signed(-13046, D_WIDTH),
        to_signed(-13300, D_WIDTH),
        to_signed(-13552, D_WIDTH),
        to_signed(-13801, D_WIDTH),
        to_signed(-14047, D_WIDTH),
        to_signed(-14290, D_WIDTH),
        to_signed(-14530, D_WIDTH),
        to_signed(-14767, D_WIDTH),
        to_signed(-15000, D_WIDTH),
        to_signed(-15230, D_WIDTH),
        to_signed(-15457, D_WIDTH),
        to_signed(-15680, D_WIDTH),
        to_signed(-15900, D_WIDTH),
        to_signed(-16115, D_WIDTH),
        to_signed(-16327, D_WIDTH),
        to_signed(-16535, D_WIDTH),
        to_signed(-16739, D_WIDTH),
        to_signed(-16938, D_WIDTH),
        to_signed(-17133, D_WIDTH),
        to_signed(-17324, D_WIDTH),
        to_signed(-17511, D_WIDTH),
        to_signed(-17693, D_WIDTH),
        to_signed(-17870, D_WIDTH),
        to_signed(-18042, D_WIDTH),
        to_signed(-18210, D_WIDTH),
        to_signed(-18373, D_WIDTH),
        to_signed(-18530, D_WIDTH),
        to_signed(-18683, D_WIDTH),
        to_signed(-18830, D_WIDTH),
        to_signed(-18972, D_WIDTH),
        to_signed(-19109, D_WIDTH),
        to_signed(-19240, D_WIDTH),
        to_signed(-19365, D_WIDTH),
        to_signed(-19485, D_WIDTH),
        to_signed(-19599, D_WIDTH),
        to_signed(-19707, D_WIDTH),
        to_signed(-19810, D_WIDTH),
        to_signed(-19906, D_WIDTH),
        to_signed(-19997, D_WIDTH),
        to_signed(-20081, D_WIDTH),
        to_signed(-20159, D_WIDTH),
        to_signed(-20230, D_WIDTH),
        to_signed(-20295, D_WIDTH),
        to_signed(-20354, D_WIDTH),
        to_signed(-20406, D_WIDTH),
        to_signed(-20452, D_WIDTH),
        to_signed(-20491, D_WIDTH),
        to_signed(-20523, D_WIDTH),
        to_signed(-20548, D_WIDTH),
        to_signed(-20566, D_WIDTH),
        to_signed(-20578, D_WIDTH),
        to_signed(-20582, D_WIDTH),
        to_signed(-20579, D_WIDTH),
        to_signed(-20570, D_WIDTH),
        to_signed(-20552, D_WIDTH),
        to_signed(-20528, D_WIDTH),
        to_signed(-20496, D_WIDTH),
        to_signed(-20457, D_WIDTH),
        to_signed(-20411, D_WIDTH),
        to_signed(-20357, D_WIDTH),
        to_signed(-20295, D_WIDTH),
        to_signed(-20226, D_WIDTH),
        to_signed(-20149, D_WIDTH),
        to_signed(-20064, D_WIDTH),
        to_signed(-19972, D_WIDTH),
        to_signed(-19872, D_WIDTH),
        to_signed(-19764, D_WIDTH),
        to_signed(-19648, D_WIDTH),
        to_signed(-19524, D_WIDTH),
        to_signed(-19392, D_WIDTH),
        to_signed(-19253, D_WIDTH),
        to_signed(-19105, D_WIDTH),
        to_signed(-18949, D_WIDTH),
        to_signed(-18786, D_WIDTH),
        to_signed(-18614, D_WIDTH),
        to_signed(-18434, D_WIDTH),
        to_signed(-18245, D_WIDTH),
        to_signed(-18049, D_WIDTH),
        to_signed(-17844, D_WIDTH),
        to_signed(-17632, D_WIDTH),
        to_signed(-17411, D_WIDTH),
        to_signed(-17181, D_WIDTH),
        to_signed(-16944, D_WIDTH),
        to_signed(-16698, D_WIDTH),
        to_signed(-16444, D_WIDTH),
        to_signed(-16181, D_WIDTH),
        to_signed(-15911, D_WIDTH),
        to_signed(-15632, D_WIDTH),
        to_signed(-15345, D_WIDTH),
        to_signed(-15049, D_WIDTH),
        to_signed(-14745, D_WIDTH),
        to_signed(-14433, D_WIDTH),
        to_signed(-14113, D_WIDTH),
        to_signed(-13784, D_WIDTH),
        to_signed(-13447, D_WIDTH),
        to_signed(-13102, D_WIDTH),
        to_signed(-12749, D_WIDTH),
        to_signed(-12387, D_WIDTH),
        to_signed(-12017, D_WIDTH),
        to_signed(-11639, D_WIDTH),
        to_signed(-11253, D_WIDTH),
        to_signed(-10859, D_WIDTH),
        to_signed(-10457, D_WIDTH),
        to_signed(-10047, D_WIDTH),
        to_signed(-9628, D_WIDTH),
        to_signed(-9202, D_WIDTH),
        to_signed(-8768, D_WIDTH),
        to_signed(-8325, D_WIDTH),
        to_signed(-7875, D_WIDTH),
        to_signed(-7417, D_WIDTH),
        to_signed(-6951, D_WIDTH),
        to_signed(-6478, D_WIDTH),
        to_signed(-5997, D_WIDTH),
        to_signed(-5508, D_WIDTH),
        to_signed(-5012, D_WIDTH),
        to_signed(-4508, D_WIDTH),
        to_signed(-3996, D_WIDTH),
        to_signed(-3477, D_WIDTH),
        to_signed(-2951, D_WIDTH),
        to_signed(-2417, D_WIDTH),
        to_signed(-1877, D_WIDTH),
        to_signed(-1329, D_WIDTH),
        to_signed(-773, D_WIDTH),
        to_signed(-211, D_WIDTH),
        to_signed(358, D_WIDTH),
        to_signed(934, D_WIDTH),
        to_signed(1517, D_WIDTH),
        to_signed(2106, D_WIDTH),
        to_signed(2702, D_WIDTH),
        to_signed(3305, D_WIDTH),
        to_signed(3914, D_WIDTH),
        to_signed(4530, D_WIDTH),
        to_signed(5152, D_WIDTH),
        to_signed(5780, D_WIDTH),
        to_signed(6415, D_WIDTH),
        to_signed(7055, D_WIDTH),
        to_signed(7701, D_WIDTH),
        to_signed(8354, D_WIDTH),
        to_signed(9012, D_WIDTH),
        to_signed(9675, D_WIDTH),
        to_signed(10344, D_WIDTH),
        to_signed(11019, D_WIDTH),
        to_signed(11699, D_WIDTH),
        to_signed(12384, D_WIDTH),
        to_signed(13075, D_WIDTH),
        to_signed(13770, D_WIDTH),
        to_signed(14471, D_WIDTH),
        to_signed(15176, D_WIDTH),
        to_signed(15886, D_WIDTH),
        to_signed(16600, D_WIDTH),
        to_signed(17319, D_WIDTH),
        to_signed(18043, D_WIDTH),
        to_signed(18770, D_WIDTH),
        to_signed(19502, D_WIDTH),
        to_signed(20237, D_WIDTH),
        to_signed(20977, D_WIDTH),
        to_signed(21720, D_WIDTH),
        to_signed(22467, D_WIDTH),
        to_signed(23217, D_WIDTH),
        to_signed(23971, D_WIDTH),
        to_signed(24728, D_WIDTH),
        to_signed(25488, D_WIDTH),
        to_signed(26251, D_WIDTH),
        to_signed(27017, D_WIDTH),
        to_signed(27785, D_WIDTH),
        to_signed(28556, D_WIDTH),
        to_signed(29330, D_WIDTH),
        to_signed(30106, D_WIDTH),
        to_signed(30884, D_WIDTH),
        to_signed(31664, D_WIDTH),
        to_signed(32446, D_WIDTH),
        to_signed(33229, D_WIDTH),
        to_signed(34015, D_WIDTH),
        to_signed(34801, D_WIDTH),
        to_signed(35589, D_WIDTH),
        to_signed(36379, D_WIDTH),
        to_signed(37169, D_WIDTH),
        to_signed(37960, D_WIDTH),
        to_signed(38752, D_WIDTH),
        to_signed(39544, D_WIDTH),
        to_signed(40337, D_WIDTH),
        to_signed(41130, D_WIDTH),
        to_signed(41923, D_WIDTH),
        to_signed(42717, D_WIDTH),
        to_signed(43510, D_WIDTH),
        to_signed(44303, D_WIDTH),
        to_signed(45095, D_WIDTH),
        to_signed(45887, D_WIDTH),
        to_signed(46678, D_WIDTH),
        to_signed(47468, D_WIDTH),
        to_signed(48257, D_WIDTH),
        to_signed(49045, D_WIDTH),
        to_signed(49832, D_WIDTH),
        to_signed(50617, D_WIDTH),
        to_signed(51400, D_WIDTH),
        to_signed(52182, D_WIDTH),
        to_signed(52962, D_WIDTH),
        to_signed(53739, D_WIDTH),
        to_signed(54515, D_WIDTH),
        to_signed(55288, D_WIDTH),
        to_signed(56058, D_WIDTH),
        to_signed(56826, D_WIDTH),
        to_signed(57591, D_WIDTH),
        to_signed(58353, D_WIDTH),
        to_signed(59111, D_WIDTH),
        to_signed(59867, D_WIDTH),
        to_signed(60619, D_WIDTH),
        to_signed(61367, D_WIDTH),
        to_signed(62112, D_WIDTH),
        to_signed(62853, D_WIDTH),
        to_signed(63589, D_WIDTH),
        to_signed(64322, D_WIDTH),
        to_signed(65050, D_WIDTH),
        to_signed(65774, D_WIDTH),
        to_signed(66493, D_WIDTH),
        to_signed(67208, D_WIDTH),
        to_signed(67917, D_WIDTH),
        to_signed(68622, D_WIDTH),
        to_signed(69321, D_WIDTH),
        to_signed(70015, D_WIDTH),
        to_signed(70703, D_WIDTH),
        to_signed(71386, D_WIDTH),
        to_signed(72063, D_WIDTH),
        to_signed(72735, D_WIDTH),
        to_signed(73400, D_WIDTH),
        to_signed(74059, D_WIDTH),
        to_signed(74712, D_WIDTH),
        to_signed(75358, D_WIDTH),
        to_signed(75998, D_WIDTH),
        to_signed(76632, D_WIDTH),
        to_signed(77258, D_WIDTH),
        to_signed(77878, D_WIDTH),
        to_signed(78490, D_WIDTH),
        to_signed(79095, D_WIDTH),
        to_signed(79693, D_WIDTH),
        to_signed(80284, D_WIDTH),
        to_signed(80867, D_WIDTH),
        to_signed(81442, D_WIDTH),
        to_signed(82010, D_WIDTH),
        to_signed(82570, D_WIDTH),
        to_signed(83121, D_WIDTH),
        to_signed(83665, D_WIDTH),
        to_signed(84200, D_WIDTH),
        to_signed(84727, D_WIDTH),
        to_signed(85246, D_WIDTH),
        to_signed(85756, D_WIDTH),
        to_signed(86257, D_WIDTH),
        to_signed(86750, D_WIDTH),
        to_signed(87233, D_WIDTH),
        to_signed(87708, D_WIDTH),
        to_signed(88174, D_WIDTH),
        to_signed(88630, D_WIDTH),
        to_signed(89077, D_WIDTH),
        to_signed(89515, D_WIDTH),
        to_signed(89943, D_WIDTH),
        to_signed(90362, D_WIDTH),
        to_signed(90772, D_WIDTH),
        to_signed(91171, D_WIDTH),
        to_signed(91561, D_WIDTH),
        to_signed(91941, D_WIDTH),
        to_signed(92311, D_WIDTH),
        to_signed(92670, D_WIDTH),
        to_signed(93020, D_WIDTH),
        to_signed(93360, D_WIDTH),
        to_signed(93689, D_WIDTH),
        to_signed(94008, D_WIDTH),
        to_signed(94317, D_WIDTH),
        to_signed(94615, D_WIDTH),
        to_signed(94903, D_WIDTH),
        to_signed(95180, D_WIDTH),
        to_signed(95446, D_WIDTH),
        to_signed(95702, D_WIDTH),
        to_signed(95947, D_WIDTH),
        to_signed(96182, D_WIDTH),
        to_signed(96405, D_WIDTH),
        to_signed(96618, D_WIDTH),
        to_signed(96819, D_WIDTH),
        to_signed(97010, D_WIDTH),
        to_signed(97190, D_WIDTH),
        to_signed(97359, D_WIDTH),
        to_signed(97516, D_WIDTH),
        to_signed(97663, D_WIDTH),
        to_signed(97798, D_WIDTH),
        to_signed(97922, D_WIDTH),
        to_signed(98035, D_WIDTH),
        to_signed(98137, D_WIDTH),
        to_signed(98227, D_WIDTH),
        to_signed(98306, D_WIDTH),
        to_signed(98374, D_WIDTH),
        to_signed(98431, D_WIDTH),
        to_signed(98476, D_WIDTH),
        to_signed(98510, D_WIDTH),
        to_signed(98533, D_WIDTH),
        to_signed(98544, D_WIDTH),
        -- 2048 - 1920 = 128 padding works
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH)
    );

begin

    process(clk)
    begin
        if rising_edge(clk) then
            if clk_en = '1' then
                data <= coeff_list(to_integer(addr));
            end if;
        end if;
    end process;

end rtl;
