library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity coeff_rom is
    generic(
        A_WIDTH : integer;
        D_WIDTH : integer
        );
    port (
        clk    : in  std_logic;
        clk_en : in  std_logic;
        addr   : in  unsigned(A_WIDTH - 1 downto 0);
        data   : out signed(D_WIDTH - 1 downto 0)
        );
end;

architecture rtl of coeff_rom is

    type t_coeff_list is array(0 to 2 ** A_WIDTH - 1) of
        signed(D_WIDTH - 1 downto 0);

    -- In GNU Octave:
    -- f1 = 16000
    -- f2 = 24000
    -- Fsimm1 = 6000000
    -- att1 = db2mag(-60)    # Seems to be ignored
    -- att2 = db2mag(-81.5)
    -- [n,Wn,beta,ftype] = kaiserord([f1 f2], [1 0],[att1 att2], Fsimm1)
    -- hc = fir1(n-1, Wn, ftype, kaiser(n, beta));
    -- hc = hc * 2^8;
    -- hc = round(hc * 2^16);
    -- save hc.txt hc;

    signal coeff_list : t_coeff_list := (
        to_signed(5, D_WIDTH),
        to_signed(6, D_WIDTH),
        to_signed(6, D_WIDTH),
        to_signed(6, D_WIDTH),
        to_signed(6, D_WIDTH),
        to_signed(6, D_WIDTH),
        to_signed(6, D_WIDTH),
        to_signed(6, D_WIDTH),
        to_signed(6, D_WIDTH),
        to_signed(6, D_WIDTH),
        to_signed(6, D_WIDTH),
        to_signed(7, D_WIDTH),
        to_signed(7, D_WIDTH),
        to_signed(7, D_WIDTH),
        to_signed(7, D_WIDTH),
        to_signed(7, D_WIDTH),
        to_signed(7, D_WIDTH),
        to_signed(7, D_WIDTH),
        to_signed(7, D_WIDTH),
        to_signed(7, D_WIDTH),
        to_signed(7, D_WIDTH),
        to_signed(7, D_WIDTH),
        to_signed(7, D_WIDTH),
        to_signed(8, D_WIDTH),
        to_signed(8, D_WIDTH),
        to_signed(8, D_WIDTH),
        to_signed(8, D_WIDTH),
        to_signed(8, D_WIDTH),
        to_signed(8, D_WIDTH),
        to_signed(8, D_WIDTH),
        to_signed(8, D_WIDTH),
        to_signed(8, D_WIDTH),
        to_signed(8, D_WIDTH),
        to_signed(8, D_WIDTH),
        to_signed(8, D_WIDTH),
        to_signed(8, D_WIDTH),
        to_signed(8, D_WIDTH),
        to_signed(8, D_WIDTH),
        to_signed(8, D_WIDTH),
        to_signed(8, D_WIDTH),
        to_signed(8, D_WIDTH),
        to_signed(8, D_WIDTH),
        to_signed(8, D_WIDTH),
        to_signed(8, D_WIDTH),
        to_signed(8, D_WIDTH),
        to_signed(8, D_WIDTH),
        to_signed(8, D_WIDTH),
        to_signed(8, D_WIDTH),
        to_signed(7, D_WIDTH),
        to_signed(7, D_WIDTH),
        to_signed(7, D_WIDTH),
        to_signed(7, D_WIDTH),
        to_signed(7, D_WIDTH),
        to_signed(7, D_WIDTH),
        to_signed(7, D_WIDTH),
        to_signed(7, D_WIDTH),
        to_signed(7, D_WIDTH),
        to_signed(6, D_WIDTH),
        to_signed(6, D_WIDTH),
        to_signed(6, D_WIDTH),
        to_signed(6, D_WIDTH),
        to_signed(6, D_WIDTH),
        to_signed(6, D_WIDTH),
        to_signed(6, D_WIDTH),
        to_signed(5, D_WIDTH),
        to_signed(5, D_WIDTH),
        to_signed(5, D_WIDTH),
        to_signed(5, D_WIDTH),
        to_signed(5, D_WIDTH),
        to_signed(4, D_WIDTH),
        to_signed(4, D_WIDTH),
        to_signed(4, D_WIDTH),
        to_signed(4, D_WIDTH),
        to_signed(3, D_WIDTH),
        to_signed(3, D_WIDTH),
        to_signed(3, D_WIDTH),
        to_signed(2, D_WIDTH),
        to_signed(2, D_WIDTH),
        to_signed(2, D_WIDTH),
        to_signed(2, D_WIDTH),
        to_signed(1, D_WIDTH),
        to_signed(1, D_WIDTH),
        to_signed(1, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(-0, D_WIDTH),
        to_signed(-0, D_WIDTH),
        to_signed(-1, D_WIDTH),
        to_signed(-1, D_WIDTH),
        to_signed(-2, D_WIDTH),
        to_signed(-2, D_WIDTH),
        to_signed(-2, D_WIDTH),
        to_signed(-3, D_WIDTH),
        to_signed(-3, D_WIDTH),
        to_signed(-4, D_WIDTH),
        to_signed(-4, D_WIDTH),
        to_signed(-4, D_WIDTH),
        to_signed(-5, D_WIDTH),
        to_signed(-5, D_WIDTH),
        to_signed(-6, D_WIDTH),
        to_signed(-6, D_WIDTH),
        to_signed(-7, D_WIDTH),
        to_signed(-7, D_WIDTH),
        to_signed(-8, D_WIDTH),
        to_signed(-8, D_WIDTH),
        to_signed(-8, D_WIDTH),
        to_signed(-9, D_WIDTH),
        to_signed(-9, D_WIDTH),
        to_signed(-10, D_WIDTH),
        to_signed(-10, D_WIDTH),
        to_signed(-11, D_WIDTH),
        to_signed(-11, D_WIDTH),
        to_signed(-12, D_WIDTH),
        to_signed(-12, D_WIDTH),
        to_signed(-13, D_WIDTH),
        to_signed(-14, D_WIDTH),
        to_signed(-14, D_WIDTH),
        to_signed(-15, D_WIDTH),
        to_signed(-15, D_WIDTH),
        to_signed(-16, D_WIDTH),
        to_signed(-16, D_WIDTH),
        to_signed(-17, D_WIDTH),
        to_signed(-17, D_WIDTH),
        to_signed(-18, D_WIDTH),
        to_signed(-18, D_WIDTH),
        to_signed(-19, D_WIDTH),
        to_signed(-19, D_WIDTH),
        to_signed(-20, D_WIDTH),
        to_signed(-20, D_WIDTH),
        to_signed(-21, D_WIDTH),
        to_signed(-21, D_WIDTH),
        to_signed(-22, D_WIDTH),
        to_signed(-23, D_WIDTH),
        to_signed(-23, D_WIDTH),
        to_signed(-24, D_WIDTH),
        to_signed(-24, D_WIDTH),
        to_signed(-25, D_WIDTH),
        to_signed(-25, D_WIDTH),
        to_signed(-26, D_WIDTH),
        to_signed(-26, D_WIDTH),
        to_signed(-27, D_WIDTH),
        to_signed(-27, D_WIDTH),
        to_signed(-28, D_WIDTH),
        to_signed(-28, D_WIDTH),
        to_signed(-29, D_WIDTH),
        to_signed(-29, D_WIDTH),
        to_signed(-30, D_WIDTH),
        to_signed(-30, D_WIDTH),
        to_signed(-30, D_WIDTH),
        to_signed(-31, D_WIDTH),
        to_signed(-31, D_WIDTH),
        to_signed(-32, D_WIDTH),
        to_signed(-32, D_WIDTH),
        to_signed(-33, D_WIDTH),
        to_signed(-33, D_WIDTH),
        to_signed(-33, D_WIDTH),
        to_signed(-34, D_WIDTH),
        to_signed(-34, D_WIDTH),
        to_signed(-34, D_WIDTH),
        to_signed(-35, D_WIDTH),
        to_signed(-35, D_WIDTH),
        to_signed(-35, D_WIDTH),
        to_signed(-36, D_WIDTH),
        to_signed(-36, D_WIDTH),
        to_signed(-36, D_WIDTH),
        to_signed(-37, D_WIDTH),
        to_signed(-37, D_WIDTH),
        to_signed(-37, D_WIDTH),
        to_signed(-37, D_WIDTH),
        to_signed(-38, D_WIDTH),
        to_signed(-38, D_WIDTH),
        to_signed(-38, D_WIDTH),
        to_signed(-38, D_WIDTH),
        to_signed(-38, D_WIDTH),
        to_signed(-38, D_WIDTH),
        to_signed(-38, D_WIDTH),
        to_signed(-38, D_WIDTH),
        to_signed(-39, D_WIDTH),
        to_signed(-39, D_WIDTH),
        to_signed(-39, D_WIDTH),
        to_signed(-39, D_WIDTH),
        to_signed(-39, D_WIDTH),
        to_signed(-39, D_WIDTH),
        to_signed(-39, D_WIDTH),
        to_signed(-38, D_WIDTH),
        to_signed(-38, D_WIDTH),
        to_signed(-38, D_WIDTH),
        to_signed(-38, D_WIDTH),
        to_signed(-38, D_WIDTH),
        to_signed(-38, D_WIDTH),
        to_signed(-38, D_WIDTH),
        to_signed(-37, D_WIDTH),
        to_signed(-37, D_WIDTH),
        to_signed(-37, D_WIDTH),
        to_signed(-37, D_WIDTH),
        to_signed(-36, D_WIDTH),
        to_signed(-36, D_WIDTH),
        to_signed(-36, D_WIDTH),
        to_signed(-35, D_WIDTH),
        to_signed(-35, D_WIDTH),
        to_signed(-34, D_WIDTH),
        to_signed(-34, D_WIDTH),
        to_signed(-33, D_WIDTH),
        to_signed(-33, D_WIDTH),
        to_signed(-32, D_WIDTH),
        to_signed(-32, D_WIDTH),
        to_signed(-31, D_WIDTH),
        to_signed(-31, D_WIDTH),
        to_signed(-30, D_WIDTH),
        to_signed(-29, D_WIDTH),
        to_signed(-29, D_WIDTH),
        to_signed(-28, D_WIDTH),
        to_signed(-27, D_WIDTH),
        to_signed(-27, D_WIDTH),
        to_signed(-26, D_WIDTH),
        to_signed(-25, D_WIDTH),
        to_signed(-24, D_WIDTH),
        to_signed(-23, D_WIDTH),
        to_signed(-22, D_WIDTH),
        to_signed(-22, D_WIDTH),
        to_signed(-21, D_WIDTH),
        to_signed(-20, D_WIDTH),
        to_signed(-19, D_WIDTH),
        to_signed(-18, D_WIDTH),
        to_signed(-17, D_WIDTH),
        to_signed(-16, D_WIDTH),
        to_signed(-15, D_WIDTH),
        to_signed(-14, D_WIDTH),
        to_signed(-12, D_WIDTH),
        to_signed(-11, D_WIDTH),
        to_signed(-10, D_WIDTH),
        to_signed(-9, D_WIDTH),
        to_signed(-8, D_WIDTH),
        to_signed(-7, D_WIDTH),
        to_signed(-5, D_WIDTH),
        to_signed(-4, D_WIDTH),
        to_signed(-3, D_WIDTH),
        to_signed(-1, D_WIDTH),
        to_signed(-0, D_WIDTH),
        to_signed(1, D_WIDTH),
        to_signed(3, D_WIDTH),
        to_signed(4, D_WIDTH),
        to_signed(5, D_WIDTH),
        to_signed(7, D_WIDTH),
        to_signed(8, D_WIDTH),
        to_signed(10, D_WIDTH),
        to_signed(11, D_WIDTH),
        to_signed(13, D_WIDTH),
        to_signed(14, D_WIDTH),
        to_signed(16, D_WIDTH),
        to_signed(17, D_WIDTH),
        to_signed(19, D_WIDTH),
        to_signed(20, D_WIDTH),
        to_signed(22, D_WIDTH),
        to_signed(23, D_WIDTH),
        to_signed(25, D_WIDTH),
        to_signed(27, D_WIDTH),
        to_signed(28, D_WIDTH),
        to_signed(30, D_WIDTH),
        to_signed(31, D_WIDTH),
        to_signed(33, D_WIDTH),
        to_signed(35, D_WIDTH),
        to_signed(36, D_WIDTH),
        to_signed(38, D_WIDTH),
        to_signed(40, D_WIDTH),
        to_signed(41, D_WIDTH),
        to_signed(43, D_WIDTH),
        to_signed(45, D_WIDTH),
        to_signed(46, D_WIDTH),
        to_signed(48, D_WIDTH),
        to_signed(50, D_WIDTH),
        to_signed(51, D_WIDTH),
        to_signed(53, D_WIDTH),
        to_signed(55, D_WIDTH),
        to_signed(56, D_WIDTH),
        to_signed(58, D_WIDTH),
        to_signed(60, D_WIDTH),
        to_signed(61, D_WIDTH),
        to_signed(63, D_WIDTH),
        to_signed(65, D_WIDTH),
        to_signed(66, D_WIDTH),
        to_signed(68, D_WIDTH),
        to_signed(69, D_WIDTH),
        to_signed(71, D_WIDTH),
        to_signed(72, D_WIDTH),
        to_signed(74, D_WIDTH),
        to_signed(76, D_WIDTH),
        to_signed(77, D_WIDTH),
        to_signed(79, D_WIDTH),
        to_signed(80, D_WIDTH),
        to_signed(82, D_WIDTH),
        to_signed(83, D_WIDTH),
        to_signed(85, D_WIDTH),
        to_signed(86, D_WIDTH),
        to_signed(87, D_WIDTH),
        to_signed(89, D_WIDTH),
        to_signed(90, D_WIDTH),
        to_signed(91, D_WIDTH),
        to_signed(93, D_WIDTH),
        to_signed(94, D_WIDTH),
        to_signed(95, D_WIDTH),
        to_signed(96, D_WIDTH),
        to_signed(98, D_WIDTH),
        to_signed(99, D_WIDTH),
        to_signed(100, D_WIDTH),
        to_signed(101, D_WIDTH),
        to_signed(102, D_WIDTH),
        to_signed(103, D_WIDTH),
        to_signed(104, D_WIDTH),
        to_signed(105, D_WIDTH),
        to_signed(106, D_WIDTH),
        to_signed(107, D_WIDTH),
        to_signed(108, D_WIDTH),
        to_signed(108, D_WIDTH),
        to_signed(109, D_WIDTH),
        to_signed(110, D_WIDTH),
        to_signed(110, D_WIDTH),
        to_signed(111, D_WIDTH),
        to_signed(112, D_WIDTH),
        to_signed(112, D_WIDTH),
        to_signed(113, D_WIDTH),
        to_signed(113, D_WIDTH),
        to_signed(113, D_WIDTH),
        to_signed(114, D_WIDTH),
        to_signed(114, D_WIDTH),
        to_signed(114, D_WIDTH),
        to_signed(115, D_WIDTH),
        to_signed(115, D_WIDTH),
        to_signed(115, D_WIDTH),
        to_signed(115, D_WIDTH),
        to_signed(115, D_WIDTH),
        to_signed(115, D_WIDTH),
        to_signed(115, D_WIDTH),
        to_signed(114, D_WIDTH),
        to_signed(114, D_WIDTH),
        to_signed(114, D_WIDTH),
        to_signed(113, D_WIDTH),
        to_signed(113, D_WIDTH),
        to_signed(113, D_WIDTH),
        to_signed(112, D_WIDTH),
        to_signed(111, D_WIDTH),
        to_signed(111, D_WIDTH),
        to_signed(110, D_WIDTH),
        to_signed(109, D_WIDTH),
        to_signed(108, D_WIDTH),
        to_signed(108, D_WIDTH),
        to_signed(107, D_WIDTH),
        to_signed(106, D_WIDTH),
        to_signed(104, D_WIDTH),
        to_signed(103, D_WIDTH),
        to_signed(102, D_WIDTH),
        to_signed(101, D_WIDTH),
        to_signed(100, D_WIDTH),
        to_signed(98, D_WIDTH),
        to_signed(97, D_WIDTH),
        to_signed(95, D_WIDTH),
        to_signed(94, D_WIDTH),
        to_signed(92, D_WIDTH),
        to_signed(90, D_WIDTH),
        to_signed(88, D_WIDTH),
        to_signed(87, D_WIDTH),
        to_signed(85, D_WIDTH),
        to_signed(83, D_WIDTH),
        to_signed(81, D_WIDTH),
        to_signed(79, D_WIDTH),
        to_signed(77, D_WIDTH),
        to_signed(74, D_WIDTH),
        to_signed(72, D_WIDTH),
        to_signed(70, D_WIDTH),
        to_signed(67, D_WIDTH),
        to_signed(65, D_WIDTH),
        to_signed(62, D_WIDTH),
        to_signed(60, D_WIDTH),
        to_signed(57, D_WIDTH),
        to_signed(55, D_WIDTH),
        to_signed(52, D_WIDTH),
        to_signed(49, D_WIDTH),
        to_signed(46, D_WIDTH),
        to_signed(43, D_WIDTH),
        to_signed(40, D_WIDTH),
        to_signed(37, D_WIDTH),
        to_signed(34, D_WIDTH),
        to_signed(31, D_WIDTH),
        to_signed(28, D_WIDTH),
        to_signed(25, D_WIDTH),
        to_signed(22, D_WIDTH),
        to_signed(18, D_WIDTH),
        to_signed(15, D_WIDTH),
        to_signed(12, D_WIDTH),
        to_signed(8, D_WIDTH),
        to_signed(5, D_WIDTH),
        to_signed(1, D_WIDTH),
        to_signed(-2, D_WIDTH),
        to_signed(-6, D_WIDTH),
        to_signed(-10, D_WIDTH),
        to_signed(-13, D_WIDTH),
        to_signed(-17, D_WIDTH),
        to_signed(-21, D_WIDTH),
        to_signed(-25, D_WIDTH),
        to_signed(-28, D_WIDTH),
        to_signed(-32, D_WIDTH),
        to_signed(-36, D_WIDTH),
        to_signed(-40, D_WIDTH),
        to_signed(-44, D_WIDTH),
        to_signed(-48, D_WIDTH),
        to_signed(-52, D_WIDTH),
        to_signed(-56, D_WIDTH),
        to_signed(-60, D_WIDTH),
        to_signed(-64, D_WIDTH),
        to_signed(-68, D_WIDTH),
        to_signed(-72, D_WIDTH),
        to_signed(-76, D_WIDTH),
        to_signed(-80, D_WIDTH),
        to_signed(-84, D_WIDTH),
        to_signed(-88, D_WIDTH),
        to_signed(-92, D_WIDTH),
        to_signed(-97, D_WIDTH),
        to_signed(-101, D_WIDTH),
        to_signed(-105, D_WIDTH),
        to_signed(-109, D_WIDTH),
        to_signed(-113, D_WIDTH),
        to_signed(-117, D_WIDTH),
        to_signed(-121, D_WIDTH),
        to_signed(-125, D_WIDTH),
        to_signed(-129, D_WIDTH),
        to_signed(-133, D_WIDTH),
        to_signed(-137, D_WIDTH),
        to_signed(-141, D_WIDTH),
        to_signed(-145, D_WIDTH),
        to_signed(-149, D_WIDTH),
        to_signed(-153, D_WIDTH),
        to_signed(-157, D_WIDTH),
        to_signed(-161, D_WIDTH),
        to_signed(-165, D_WIDTH),
        to_signed(-169, D_WIDTH),
        to_signed(-172, D_WIDTH),
        to_signed(-176, D_WIDTH),
        to_signed(-180, D_WIDTH),
        to_signed(-184, D_WIDTH),
        to_signed(-187, D_WIDTH),
        to_signed(-191, D_WIDTH),
        to_signed(-194, D_WIDTH),
        to_signed(-198, D_WIDTH),
        to_signed(-201, D_WIDTH),
        to_signed(-204, D_WIDTH),
        to_signed(-208, D_WIDTH),
        to_signed(-211, D_WIDTH),
        to_signed(-214, D_WIDTH),
        to_signed(-217, D_WIDTH),
        to_signed(-220, D_WIDTH),
        to_signed(-223, D_WIDTH),
        to_signed(-226, D_WIDTH),
        to_signed(-229, D_WIDTH),
        to_signed(-232, D_WIDTH),
        to_signed(-234, D_WIDTH),
        to_signed(-237, D_WIDTH),
        to_signed(-240, D_WIDTH),
        to_signed(-242, D_WIDTH),
        to_signed(-244, D_WIDTH),
        to_signed(-247, D_WIDTH),
        to_signed(-249, D_WIDTH),
        to_signed(-251, D_WIDTH),
        to_signed(-253, D_WIDTH),
        to_signed(-255, D_WIDTH),
        to_signed(-257, D_WIDTH),
        to_signed(-258, D_WIDTH),
        to_signed(-260, D_WIDTH),
        to_signed(-261, D_WIDTH),
        to_signed(-263, D_WIDTH),
        to_signed(-264, D_WIDTH),
        to_signed(-265, D_WIDTH),
        to_signed(-266, D_WIDTH),
        to_signed(-267, D_WIDTH),
        to_signed(-268, D_WIDTH),
        to_signed(-269, D_WIDTH),
        to_signed(-269, D_WIDTH),
        to_signed(-270, D_WIDTH),
        to_signed(-270, D_WIDTH),
        to_signed(-271, D_WIDTH),
        to_signed(-271, D_WIDTH),
        to_signed(-271, D_WIDTH),
        to_signed(-271, D_WIDTH),
        to_signed(-271, D_WIDTH),
        to_signed(-270, D_WIDTH),
        to_signed(-270, D_WIDTH),
        to_signed(-269, D_WIDTH),
        to_signed(-268, D_WIDTH),
        to_signed(-268, D_WIDTH),
        to_signed(-267, D_WIDTH),
        to_signed(-265, D_WIDTH),
        to_signed(-264, D_WIDTH),
        to_signed(-263, D_WIDTH),
        to_signed(-261, D_WIDTH),
        to_signed(-260, D_WIDTH),
        to_signed(-258, D_WIDTH),
        to_signed(-256, D_WIDTH),
        to_signed(-254, D_WIDTH),
        to_signed(-252, D_WIDTH),
        to_signed(-249, D_WIDTH),
        to_signed(-247, D_WIDTH),
        to_signed(-244, D_WIDTH),
        to_signed(-242, D_WIDTH),
        to_signed(-239, D_WIDTH),
        to_signed(-236, D_WIDTH),
        to_signed(-233, D_WIDTH),
        to_signed(-229, D_WIDTH),
        to_signed(-226, D_WIDTH),
        to_signed(-222, D_WIDTH),
        to_signed(-219, D_WIDTH),
        to_signed(-215, D_WIDTH),
        to_signed(-211, D_WIDTH),
        to_signed(-207, D_WIDTH),
        to_signed(-203, D_WIDTH),
        to_signed(-198, D_WIDTH),
        to_signed(-194, D_WIDTH),
        to_signed(-189, D_WIDTH),
        to_signed(-184, D_WIDTH),
        to_signed(-179, D_WIDTH),
        to_signed(-174, D_WIDTH),
        to_signed(-169, D_WIDTH),
        to_signed(-164, D_WIDTH),
        to_signed(-159, D_WIDTH),
        to_signed(-153, D_WIDTH),
        to_signed(-147, D_WIDTH),
        to_signed(-142, D_WIDTH),
        to_signed(-136, D_WIDTH),
        to_signed(-130, D_WIDTH),
        to_signed(-124, D_WIDTH),
        to_signed(-117, D_WIDTH),
        to_signed(-111, D_WIDTH),
        to_signed(-105, D_WIDTH),
        to_signed(-98, D_WIDTH),
        to_signed(-91, D_WIDTH),
        to_signed(-85, D_WIDTH),
        to_signed(-78, D_WIDTH),
        to_signed(-71, D_WIDTH),
        to_signed(-64, D_WIDTH),
        to_signed(-56, D_WIDTH),
        to_signed(-49, D_WIDTH),
        to_signed(-42, D_WIDTH),
        to_signed(-34, D_WIDTH),
        to_signed(-27, D_WIDTH),
        to_signed(-19, D_WIDTH),
        to_signed(-11, D_WIDTH),
        to_signed(-4, D_WIDTH),
        to_signed(4, D_WIDTH),
        to_signed(12, D_WIDTH),
        to_signed(20, D_WIDTH),
        to_signed(28, D_WIDTH),
        to_signed(36, D_WIDTH),
        to_signed(45, D_WIDTH),
        to_signed(53, D_WIDTH),
        to_signed(61, D_WIDTH),
        to_signed(70, D_WIDTH),
        to_signed(78, D_WIDTH),
        to_signed(86, D_WIDTH),
        to_signed(95, D_WIDTH),
        to_signed(103, D_WIDTH),
        to_signed(112, D_WIDTH),
        to_signed(121, D_WIDTH),
        to_signed(129, D_WIDTH),
        to_signed(138, D_WIDTH),
        to_signed(147, D_WIDTH),
        to_signed(155, D_WIDTH),
        to_signed(164, D_WIDTH),
        to_signed(173, D_WIDTH),
        to_signed(181, D_WIDTH),
        to_signed(190, D_WIDTH),
        to_signed(199, D_WIDTH),
        to_signed(207, D_WIDTH),
        to_signed(216, D_WIDTH),
        to_signed(225, D_WIDTH),
        to_signed(233, D_WIDTH),
        to_signed(242, D_WIDTH),
        to_signed(251, D_WIDTH),
        to_signed(259, D_WIDTH),
        to_signed(268, D_WIDTH),
        to_signed(276, D_WIDTH),
        to_signed(284, D_WIDTH),
        to_signed(293, D_WIDTH),
        to_signed(301, D_WIDTH),
        to_signed(309, D_WIDTH),
        to_signed(318, D_WIDTH),
        to_signed(326, D_WIDTH),
        to_signed(334, D_WIDTH),
        to_signed(342, D_WIDTH),
        to_signed(350, D_WIDTH),
        to_signed(357, D_WIDTH),
        to_signed(365, D_WIDTH),
        to_signed(373, D_WIDTH),
        to_signed(380, D_WIDTH),
        to_signed(388, D_WIDTH),
        to_signed(395, D_WIDTH),
        to_signed(402, D_WIDTH),
        to_signed(409, D_WIDTH),
        to_signed(416, D_WIDTH),
        to_signed(423, D_WIDTH),
        to_signed(430, D_WIDTH),
        to_signed(437, D_WIDTH),
        to_signed(443, D_WIDTH),
        to_signed(449, D_WIDTH),
        to_signed(456, D_WIDTH),
        to_signed(462, D_WIDTH),
        to_signed(467, D_WIDTH),
        to_signed(473, D_WIDTH),
        to_signed(479, D_WIDTH),
        to_signed(484, D_WIDTH),
        to_signed(489, D_WIDTH),
        to_signed(494, D_WIDTH),
        to_signed(499, D_WIDTH),
        to_signed(504, D_WIDTH),
        to_signed(509, D_WIDTH),
        to_signed(513, D_WIDTH),
        to_signed(517, D_WIDTH),
        to_signed(521, D_WIDTH),
        to_signed(525, D_WIDTH),
        to_signed(528, D_WIDTH),
        to_signed(532, D_WIDTH),
        to_signed(535, D_WIDTH),
        to_signed(538, D_WIDTH),
        to_signed(540, D_WIDTH),
        to_signed(543, D_WIDTH),
        to_signed(545, D_WIDTH),
        to_signed(547, D_WIDTH),
        to_signed(549, D_WIDTH),
        to_signed(550, D_WIDTH),
        to_signed(552, D_WIDTH),
        to_signed(553, D_WIDTH),
        to_signed(554, D_WIDTH),
        to_signed(554, D_WIDTH),
        to_signed(555, D_WIDTH),
        to_signed(555, D_WIDTH),
        to_signed(555, D_WIDTH),
        to_signed(555, D_WIDTH),
        to_signed(554, D_WIDTH),
        to_signed(553, D_WIDTH),
        to_signed(552, D_WIDTH),
        to_signed(551, D_WIDTH),
        to_signed(549, D_WIDTH),
        to_signed(547, D_WIDTH),
        to_signed(545, D_WIDTH),
        to_signed(543, D_WIDTH),
        to_signed(540, D_WIDTH),
        to_signed(537, D_WIDTH),
        to_signed(534, D_WIDTH),
        to_signed(531, D_WIDTH),
        to_signed(527, D_WIDTH),
        to_signed(523, D_WIDTH),
        to_signed(519, D_WIDTH),
        to_signed(514, D_WIDTH),
        to_signed(509, D_WIDTH),
        to_signed(504, D_WIDTH),
        to_signed(499, D_WIDTH),
        to_signed(493, D_WIDTH),
        to_signed(488, D_WIDTH),
        to_signed(481, D_WIDTH),
        to_signed(475, D_WIDTH),
        to_signed(468, D_WIDTH),
        to_signed(462, D_WIDTH),
        to_signed(454, D_WIDTH),
        to_signed(447, D_WIDTH),
        to_signed(439, D_WIDTH),
        to_signed(431, D_WIDTH),
        to_signed(423, D_WIDTH),
        to_signed(415, D_WIDTH),
        to_signed(406, D_WIDTH),
        to_signed(397, D_WIDTH),
        to_signed(388, D_WIDTH),
        to_signed(378, D_WIDTH),
        to_signed(368, D_WIDTH),
        to_signed(358, D_WIDTH),
        to_signed(348, D_WIDTH),
        to_signed(338, D_WIDTH),
        to_signed(327, D_WIDTH),
        to_signed(316, D_WIDTH),
        to_signed(305, D_WIDTH),
        to_signed(294, D_WIDTH),
        to_signed(282, D_WIDTH),
        to_signed(270, D_WIDTH),
        to_signed(258, D_WIDTH),
        to_signed(246, D_WIDTH),
        to_signed(233, D_WIDTH),
        to_signed(220, D_WIDTH),
        to_signed(208, D_WIDTH),
        to_signed(194, D_WIDTH),
        to_signed(181, D_WIDTH),
        to_signed(168, D_WIDTH),
        to_signed(154, D_WIDTH),
        to_signed(140, D_WIDTH),
        to_signed(126, D_WIDTH),
        to_signed(112, D_WIDTH),
        to_signed(98, D_WIDTH),
        to_signed(83, D_WIDTH),
        to_signed(68, D_WIDTH),
        to_signed(53, D_WIDTH),
        to_signed(38, D_WIDTH),
        to_signed(23, D_WIDTH),
        to_signed(8, D_WIDTH),
        to_signed(-7, D_WIDTH),
        to_signed(-23, D_WIDTH),
        to_signed(-38, D_WIDTH),
        to_signed(-54, D_WIDTH),
        to_signed(-70, D_WIDTH),
        to_signed(-86, D_WIDTH),
        to_signed(-102, D_WIDTH),
        to_signed(-118, D_WIDTH),
        to_signed(-134, D_WIDTH),
        to_signed(-151, D_WIDTH),
        to_signed(-167, D_WIDTH),
        to_signed(-183, D_WIDTH),
        to_signed(-200, D_WIDTH),
        to_signed(-216, D_WIDTH),
        to_signed(-233, D_WIDTH),
        to_signed(-249, D_WIDTH),
        to_signed(-266, D_WIDTH),
        to_signed(-283, D_WIDTH),
        to_signed(-299, D_WIDTH),
        to_signed(-316, D_WIDTH),
        to_signed(-332, D_WIDTH),
        to_signed(-349, D_WIDTH),
        to_signed(-366, D_WIDTH),
        to_signed(-382, D_WIDTH),
        to_signed(-399, D_WIDTH),
        to_signed(-415, D_WIDTH),
        to_signed(-431, D_WIDTH),
        to_signed(-448, D_WIDTH),
        to_signed(-464, D_WIDTH),
        to_signed(-480, D_WIDTH),
        to_signed(-496, D_WIDTH),
        to_signed(-512, D_WIDTH),
        to_signed(-528, D_WIDTH),
        to_signed(-544, D_WIDTH),
        to_signed(-560, D_WIDTH),
        to_signed(-575, D_WIDTH),
        to_signed(-591, D_WIDTH),
        to_signed(-606, D_WIDTH),
        to_signed(-621, D_WIDTH),
        to_signed(-636, D_WIDTH),
        to_signed(-651, D_WIDTH),
        to_signed(-666, D_WIDTH),
        to_signed(-680, D_WIDTH),
        to_signed(-695, D_WIDTH),
        to_signed(-709, D_WIDTH),
        to_signed(-723, D_WIDTH),
        to_signed(-737, D_WIDTH),
        to_signed(-750, D_WIDTH),
        to_signed(-763, D_WIDTH),
        to_signed(-776, D_WIDTH),
        to_signed(-789, D_WIDTH),
        to_signed(-802, D_WIDTH),
        to_signed(-814, D_WIDTH),
        to_signed(-826, D_WIDTH),
        to_signed(-838, D_WIDTH),
        to_signed(-849, D_WIDTH),
        to_signed(-861, D_WIDTH),
        to_signed(-871, D_WIDTH),
        to_signed(-882, D_WIDTH),
        to_signed(-892, D_WIDTH),
        to_signed(-902, D_WIDTH),
        to_signed(-912, D_WIDTH),
        to_signed(-921, D_WIDTH),
        to_signed(-930, D_WIDTH),
        to_signed(-939, D_WIDTH),
        to_signed(-947, D_WIDTH),
        to_signed(-955, D_WIDTH),
        to_signed(-963, D_WIDTH),
        to_signed(-970, D_WIDTH),
        to_signed(-977, D_WIDTH),
        to_signed(-983, D_WIDTH),
        to_signed(-990, D_WIDTH),
        to_signed(-995, D_WIDTH),
        to_signed(-1001, D_WIDTH),
        to_signed(-1005, D_WIDTH),
        to_signed(-1010, D_WIDTH),
        to_signed(-1014, D_WIDTH),
        to_signed(-1018, D_WIDTH),
        to_signed(-1021, D_WIDTH),
        to_signed(-1024, D_WIDTH),
        to_signed(-1026, D_WIDTH),
        to_signed(-1028, D_WIDTH),
        to_signed(-1030, D_WIDTH),
        to_signed(-1031, D_WIDTH),
        to_signed(-1031, D_WIDTH),
        to_signed(-1032, D_WIDTH),
        to_signed(-1031, D_WIDTH),
        to_signed(-1031, D_WIDTH),
        to_signed(-1030, D_WIDTH),
        to_signed(-1028, D_WIDTH),
        to_signed(-1026, D_WIDTH),
        to_signed(-1023, D_WIDTH),
        to_signed(-1020, D_WIDTH),
        to_signed(-1017, D_WIDTH),
        to_signed(-1013, D_WIDTH),
        to_signed(-1008, D_WIDTH),
        to_signed(-1003, D_WIDTH),
        to_signed(-998, D_WIDTH),
        to_signed(-992, D_WIDTH),
        to_signed(-986, D_WIDTH),
        to_signed(-979, D_WIDTH),
        to_signed(-971, D_WIDTH),
        to_signed(-964, D_WIDTH),
        to_signed(-955, D_WIDTH),
        to_signed(-946, D_WIDTH),
        to_signed(-937, D_WIDTH),
        to_signed(-927, D_WIDTH),
        to_signed(-917, D_WIDTH),
        to_signed(-906, D_WIDTH),
        to_signed(-895, D_WIDTH),
        to_signed(-884, D_WIDTH),
        to_signed(-871, D_WIDTH),
        to_signed(-859, D_WIDTH),
        to_signed(-846, D_WIDTH),
        to_signed(-832, D_WIDTH),
        to_signed(-818, D_WIDTH),
        to_signed(-804, D_WIDTH),
        to_signed(-789, D_WIDTH),
        to_signed(-773, D_WIDTH),
        to_signed(-757, D_WIDTH),
        to_signed(-741, D_WIDTH),
        to_signed(-724, D_WIDTH),
        to_signed(-707, D_WIDTH),
        to_signed(-689, D_WIDTH),
        to_signed(-671, D_WIDTH),
        to_signed(-653, D_WIDTH),
        to_signed(-634, D_WIDTH),
        to_signed(-614, D_WIDTH),
        to_signed(-595, D_WIDTH),
        to_signed(-575, D_WIDTH),
        to_signed(-554, D_WIDTH),
        to_signed(-533, D_WIDTH),
        to_signed(-512, D_WIDTH),
        to_signed(-490, D_WIDTH),
        to_signed(-468, D_WIDTH),
        to_signed(-445, D_WIDTH),
        to_signed(-422, D_WIDTH),
        to_signed(-399, D_WIDTH),
        to_signed(-376, D_WIDTH),
        to_signed(-352, D_WIDTH),
        to_signed(-328, D_WIDTH),
        to_signed(-303, D_WIDTH),
        to_signed(-278, D_WIDTH),
        to_signed(-253, D_WIDTH),
        to_signed(-228, D_WIDTH),
        to_signed(-202, D_WIDTH),
        to_signed(-176, D_WIDTH),
        to_signed(-150, D_WIDTH),
        to_signed(-123, D_WIDTH),
        to_signed(-96, D_WIDTH),
        to_signed(-69, D_WIDTH),
        to_signed(-42, D_WIDTH),
        to_signed(-15, D_WIDTH),
        to_signed(13, D_WIDTH),
        to_signed(41, D_WIDTH),
        to_signed(69, D_WIDTH),
        to_signed(97, D_WIDTH),
        to_signed(126, D_WIDTH),
        to_signed(154, D_WIDTH),
        to_signed(183, D_WIDTH),
        to_signed(212, D_WIDTH),
        to_signed(240, D_WIDTH),
        to_signed(269, D_WIDTH),
        to_signed(299, D_WIDTH),
        to_signed(328, D_WIDTH),
        to_signed(357, D_WIDTH),
        to_signed(386, D_WIDTH),
        to_signed(416, D_WIDTH),
        to_signed(445, D_WIDTH),
        to_signed(474, D_WIDTH),
        to_signed(504, D_WIDTH),
        to_signed(533, D_WIDTH),
        to_signed(562, D_WIDTH),
        to_signed(592, D_WIDTH),
        to_signed(621, D_WIDTH),
        to_signed(650, D_WIDTH),
        to_signed(679, D_WIDTH),
        to_signed(708, D_WIDTH),
        to_signed(737, D_WIDTH),
        to_signed(766, D_WIDTH),
        to_signed(795, D_WIDTH),
        to_signed(823, D_WIDTH),
        to_signed(852, D_WIDTH),
        to_signed(880, D_WIDTH),
        to_signed(908, D_WIDTH),
        to_signed(936, D_WIDTH),
        to_signed(963, D_WIDTH),
        to_signed(991, D_WIDTH),
        to_signed(1018, D_WIDTH),
        to_signed(1045, D_WIDTH),
        to_signed(1071, D_WIDTH),
        to_signed(1097, D_WIDTH),
        to_signed(1123, D_WIDTH),
        to_signed(1149, D_WIDTH),
        to_signed(1175, D_WIDTH),
        to_signed(1200, D_WIDTH),
        to_signed(1224, D_WIDTH),
        to_signed(1249, D_WIDTH),
        to_signed(1273, D_WIDTH),
        to_signed(1296, D_WIDTH),
        to_signed(1319, D_WIDTH),
        to_signed(1342, D_WIDTH),
        to_signed(1365, D_WIDTH),
        to_signed(1386, D_WIDTH),
        to_signed(1408, D_WIDTH),
        to_signed(1429, D_WIDTH),
        to_signed(1449, D_WIDTH),
        to_signed(1469, D_WIDTH),
        to_signed(1489, D_WIDTH),
        to_signed(1508, D_WIDTH),
        to_signed(1526, D_WIDTH),
        to_signed(1544, D_WIDTH),
        to_signed(1562, D_WIDTH),
        to_signed(1578, D_WIDTH),
        to_signed(1595, D_WIDTH),
        to_signed(1610, D_WIDTH),
        to_signed(1625, D_WIDTH),
        to_signed(1640, D_WIDTH),
        to_signed(1654, D_WIDTH),
        to_signed(1667, D_WIDTH),
        to_signed(1679, D_WIDTH),
        to_signed(1691, D_WIDTH),
        to_signed(1702, D_WIDTH),
        to_signed(1713, D_WIDTH),
        to_signed(1723, D_WIDTH),
        to_signed(1732, D_WIDTH),
        to_signed(1741, D_WIDTH),
        to_signed(1748, D_WIDTH),
        to_signed(1756, D_WIDTH),
        to_signed(1762, D_WIDTH),
        to_signed(1768, D_WIDTH),
        to_signed(1773, D_WIDTH),
        to_signed(1777, D_WIDTH),
        to_signed(1780, D_WIDTH),
        to_signed(1783, D_WIDTH),
        to_signed(1785, D_WIDTH),
        to_signed(1786, D_WIDTH),
        to_signed(1786, D_WIDTH),
        to_signed(1786, D_WIDTH),
        to_signed(1785, D_WIDTH),
        to_signed(1783, D_WIDTH),
        to_signed(1780, D_WIDTH),
        to_signed(1777, D_WIDTH),
        to_signed(1772, D_WIDTH),
        to_signed(1767, D_WIDTH),
        to_signed(1761, D_WIDTH),
        to_signed(1754, D_WIDTH),
        to_signed(1747, D_WIDTH),
        to_signed(1738, D_WIDTH),
        to_signed(1729, D_WIDTH),
        to_signed(1719, D_WIDTH),
        to_signed(1708, D_WIDTH),
        to_signed(1697, D_WIDTH),
        to_signed(1684, D_WIDTH),
        to_signed(1671, D_WIDTH),
        to_signed(1657, D_WIDTH),
        to_signed(1642, D_WIDTH),
        to_signed(1626, D_WIDTH),
        to_signed(1609, D_WIDTH),
        to_signed(1592, D_WIDTH),
        to_signed(1574, D_WIDTH),
        to_signed(1555, D_WIDTH),
        to_signed(1535, D_WIDTH),
        to_signed(1514, D_WIDTH),
        to_signed(1493, D_WIDTH),
        to_signed(1471, D_WIDTH),
        to_signed(1447, D_WIDTH),
        to_signed(1424, D_WIDTH),
        to_signed(1399, D_WIDTH),
        to_signed(1374, D_WIDTH),
        to_signed(1348, D_WIDTH),
        to_signed(1321, D_WIDTH),
        to_signed(1293, D_WIDTH),
        to_signed(1265, D_WIDTH),
        to_signed(1235, D_WIDTH),
        to_signed(1206, D_WIDTH),
        to_signed(1175, D_WIDTH),
        to_signed(1144, D_WIDTH),
        to_signed(1112, D_WIDTH),
        to_signed(1079, D_WIDTH),
        to_signed(1045, D_WIDTH),
        to_signed(1011, D_WIDTH),
        to_signed(977, D_WIDTH),
        to_signed(941, D_WIDTH),
        to_signed(905, D_WIDTH),
        to_signed(868, D_WIDTH),
        to_signed(831, D_WIDTH),
        to_signed(793, D_WIDTH),
        to_signed(755, D_WIDTH),
        to_signed(715, D_WIDTH),
        to_signed(676, D_WIDTH),
        to_signed(636, D_WIDTH),
        to_signed(595, D_WIDTH),
        to_signed(553, D_WIDTH),
        to_signed(512, D_WIDTH),
        to_signed(469, D_WIDTH),
        to_signed(426, D_WIDTH),
        to_signed(383, D_WIDTH),
        to_signed(339, D_WIDTH),
        to_signed(295, D_WIDTH),
        to_signed(251, D_WIDTH),
        to_signed(206, D_WIDTH),
        to_signed(160, D_WIDTH),
        to_signed(115, D_WIDTH),
        to_signed(68, D_WIDTH),
        to_signed(22, D_WIDTH),
        to_signed(-25, D_WIDTH),
        to_signed(-72, D_WIDTH),
        to_signed(-119, D_WIDTH),
        to_signed(-167, D_WIDTH),
        to_signed(-214, D_WIDTH),
        to_signed(-263, D_WIDTH),
        to_signed(-311, D_WIDTH),
        to_signed(-359, D_WIDTH),
        to_signed(-408, D_WIDTH),
        to_signed(-456, D_WIDTH),
        to_signed(-505, D_WIDTH),
        to_signed(-554, D_WIDTH),
        to_signed(-603, D_WIDTH),
        to_signed(-652, D_WIDTH),
        to_signed(-701, D_WIDTH),
        to_signed(-750, D_WIDTH),
        to_signed(-800, D_WIDTH),
        to_signed(-849, D_WIDTH),
        to_signed(-898, D_WIDTH),
        to_signed(-947, D_WIDTH),
        to_signed(-995, D_WIDTH),
        to_signed(-1044, D_WIDTH),
        to_signed(-1093, D_WIDTH),
        to_signed(-1141, D_WIDTH),
        to_signed(-1190, D_WIDTH),
        to_signed(-1238, D_WIDTH),
        to_signed(-1285, D_WIDTH),
        to_signed(-1333, D_WIDTH),
        to_signed(-1380, D_WIDTH),
        to_signed(-1427, D_WIDTH),
        to_signed(-1474, D_WIDTH),
        to_signed(-1520, D_WIDTH),
        to_signed(-1566, D_WIDTH),
        to_signed(-1612, D_WIDTH),
        to_signed(-1657, D_WIDTH),
        to_signed(-1702, D_WIDTH),
        to_signed(-1746, D_WIDTH),
        to_signed(-1790, D_WIDTH),
        to_signed(-1833, D_WIDTH),
        to_signed(-1876, D_WIDTH),
        to_signed(-1918, D_WIDTH),
        to_signed(-1960, D_WIDTH),
        to_signed(-2001, D_WIDTH),
        to_signed(-2042, D_WIDTH),
        to_signed(-2082, D_WIDTH),
        to_signed(-2121, D_WIDTH),
        to_signed(-2159, D_WIDTH),
        to_signed(-2197, D_WIDTH),
        to_signed(-2234, D_WIDTH),
        to_signed(-2271, D_WIDTH),
        to_signed(-2306, D_WIDTH),
        to_signed(-2341, D_WIDTH),
        to_signed(-2375, D_WIDTH),
        to_signed(-2409, D_WIDTH),
        to_signed(-2441, D_WIDTH),
        to_signed(-2473, D_WIDTH),
        to_signed(-2503, D_WIDTH),
        to_signed(-2533, D_WIDTH),
        to_signed(-2562, D_WIDTH),
        to_signed(-2590, D_WIDTH),
        to_signed(-2617, D_WIDTH),
        to_signed(-2643, D_WIDTH),
        to_signed(-2668, D_WIDTH),
        to_signed(-2692, D_WIDTH),
        to_signed(-2715, D_WIDTH),
        to_signed(-2737, D_WIDTH),
        to_signed(-2758, D_WIDTH),
        to_signed(-2778, D_WIDTH),
        to_signed(-2797, D_WIDTH),
        to_signed(-2815, D_WIDTH),
        to_signed(-2831, D_WIDTH),
        to_signed(-2847, D_WIDTH),
        to_signed(-2861, D_WIDTH),
        to_signed(-2874, D_WIDTH),
        to_signed(-2886, D_WIDTH),
        to_signed(-2897, D_WIDTH),
        to_signed(-2907, D_WIDTH),
        to_signed(-2915, D_WIDTH),
        to_signed(-2923, D_WIDTH),
        to_signed(-2929, D_WIDTH),
        to_signed(-2933, D_WIDTH),
        to_signed(-2937, D_WIDTH),
        to_signed(-2939, D_WIDTH),
        to_signed(-2940, D_WIDTH),
        to_signed(-2940, D_WIDTH),
        to_signed(-2938, D_WIDTH),
        to_signed(-2936, D_WIDTH),
        to_signed(-2932, D_WIDTH),
        to_signed(-2926, D_WIDTH),
        to_signed(-2919, D_WIDTH),
        to_signed(-2911, D_WIDTH),
        to_signed(-2902, D_WIDTH),
        to_signed(-2891, D_WIDTH),
        to_signed(-2879, D_WIDTH),
        to_signed(-2866, D_WIDTH),
        to_signed(-2851, D_WIDTH),
        to_signed(-2835, D_WIDTH),
        to_signed(-2818, D_WIDTH),
        to_signed(-2799, D_WIDTH),
        to_signed(-2779, D_WIDTH),
        to_signed(-2758, D_WIDTH),
        to_signed(-2735, D_WIDTH),
        to_signed(-2711, D_WIDTH),
        to_signed(-2686, D_WIDTH),
        to_signed(-2659, D_WIDTH),
        to_signed(-2632, D_WIDTH),
        to_signed(-2602, D_WIDTH),
        to_signed(-2572, D_WIDTH),
        to_signed(-2540, D_WIDTH),
        to_signed(-2507, D_WIDTH),
        to_signed(-2472, D_WIDTH),
        to_signed(-2436, D_WIDTH),
        to_signed(-2399, D_WIDTH),
        to_signed(-2361, D_WIDTH),
        to_signed(-2321, D_WIDTH),
        to_signed(-2281, D_WIDTH),
        to_signed(-2238, D_WIDTH),
        to_signed(-2195, D_WIDTH),
        to_signed(-2151, D_WIDTH),
        to_signed(-2105, D_WIDTH),
        to_signed(-2058, D_WIDTH),
        to_signed(-2010, D_WIDTH),
        to_signed(-1960, D_WIDTH),
        to_signed(-1910, D_WIDTH),
        to_signed(-1858, D_WIDTH),
        to_signed(-1806, D_WIDTH),
        to_signed(-1752, D_WIDTH),
        to_signed(-1697, D_WIDTH),
        to_signed(-1641, D_WIDTH),
        to_signed(-1584, D_WIDTH),
        to_signed(-1526, D_WIDTH),
        to_signed(-1467, D_WIDTH),
        to_signed(-1406, D_WIDTH),
        to_signed(-1345, D_WIDTH),
        to_signed(-1283, D_WIDTH),
        to_signed(-1220, D_WIDTH),
        to_signed(-1156, D_WIDTH),
        to_signed(-1091, D_WIDTH),
        to_signed(-1026, D_WIDTH),
        to_signed(-959, D_WIDTH),
        to_signed(-892, D_WIDTH),
        to_signed(-824, D_WIDTH),
        to_signed(-755, D_WIDTH),
        to_signed(-685, D_WIDTH),
        to_signed(-615, D_WIDTH),
        to_signed(-543, D_WIDTH),
        to_signed(-472, D_WIDTH),
        to_signed(-399, D_WIDTH),
        to_signed(-326, D_WIDTH),
        to_signed(-252, D_WIDTH),
        to_signed(-178, D_WIDTH),
        to_signed(-103, D_WIDTH),
        to_signed(-28, D_WIDTH),
        to_signed(48, D_WIDTH),
        to_signed(124, D_WIDTH),
        to_signed(200, D_WIDTH),
        to_signed(277, D_WIDTH),
        to_signed(355, D_WIDTH),
        to_signed(432, D_WIDTH),
        to_signed(510, D_WIDTH),
        to_signed(588, D_WIDTH),
        to_signed(667, D_WIDTH),
        to_signed(745, D_WIDTH),
        to_signed(824, D_WIDTH),
        to_signed(903, D_WIDTH),
        to_signed(982, D_WIDTH),
        to_signed(1061, D_WIDTH),
        to_signed(1140, D_WIDTH),
        to_signed(1219, D_WIDTH),
        to_signed(1298, D_WIDTH),
        to_signed(1377, D_WIDTH),
        to_signed(1456, D_WIDTH),
        to_signed(1534, D_WIDTH),
        to_signed(1613, D_WIDTH),
        to_signed(1691, D_WIDTH),
        to_signed(1769, D_WIDTH),
        to_signed(1847, D_WIDTH),
        to_signed(1924, D_WIDTH),
        to_signed(2001, D_WIDTH),
        to_signed(2077, D_WIDTH),
        to_signed(2154, D_WIDTH),
        to_signed(2229, D_WIDTH),
        to_signed(2304, D_WIDTH),
        to_signed(2379, D_WIDTH),
        to_signed(2453, D_WIDTH),
        to_signed(2527, D_WIDTH),
        to_signed(2599, D_WIDTH),
        to_signed(2672, D_WIDTH),
        to_signed(2743, D_WIDTH),
        to_signed(2814, D_WIDTH),
        to_signed(2883, D_WIDTH),
        to_signed(2952, D_WIDTH),
        to_signed(3021, D_WIDTH),
        to_signed(3088, D_WIDTH),
        to_signed(3154, D_WIDTH),
        to_signed(3219, D_WIDTH),
        to_signed(3284, D_WIDTH),
        to_signed(3347, D_WIDTH),
        to_signed(3409, D_WIDTH),
        to_signed(3471, D_WIDTH),
        to_signed(3531, D_WIDTH),
        to_signed(3589, D_WIDTH),
        to_signed(3647, D_WIDTH),
        to_signed(3703, D_WIDTH),
        to_signed(3759, D_WIDTH),
        to_signed(3813, D_WIDTH),
        to_signed(3865, D_WIDTH),
        to_signed(3916, D_WIDTH),
        to_signed(3966, D_WIDTH),
        to_signed(4014, D_WIDTH),
        to_signed(4061, D_WIDTH),
        to_signed(4107, D_WIDTH),
        to_signed(4151, D_WIDTH),
        to_signed(4193, D_WIDTH),
        to_signed(4234, D_WIDTH),
        to_signed(4273, D_WIDTH),
        to_signed(4311, D_WIDTH),
        to_signed(4347, D_WIDTH),
        to_signed(4381, D_WIDTH),
        to_signed(4414, D_WIDTH),
        to_signed(4445, D_WIDTH),
        to_signed(4474, D_WIDTH),
        to_signed(4502, D_WIDTH),
        to_signed(4527, D_WIDTH),
        to_signed(4551, D_WIDTH),
        to_signed(4573, D_WIDTH),
        to_signed(4593, D_WIDTH),
        to_signed(4612, D_WIDTH),
        to_signed(4628, D_WIDTH),
        to_signed(4642, D_WIDTH),
        to_signed(4655, D_WIDTH),
        to_signed(4666, D_WIDTH),
        to_signed(4674, D_WIDTH),
        to_signed(4681, D_WIDTH),
        to_signed(4686, D_WIDTH),
        to_signed(4689, D_WIDTH),
        to_signed(4689, D_WIDTH),
        to_signed(4688, D_WIDTH),
        to_signed(4685, D_WIDTH),
        to_signed(4679, D_WIDTH),
        to_signed(4672, D_WIDTH),
        to_signed(4662, D_WIDTH),
        to_signed(4651, D_WIDTH),
        to_signed(4637, D_WIDTH),
        to_signed(4621, D_WIDTH),
        to_signed(4603, D_WIDTH),
        to_signed(4583, D_WIDTH),
        to_signed(4561, D_WIDTH),
        to_signed(4537, D_WIDTH),
        to_signed(4511, D_WIDTH),
        to_signed(4482, D_WIDTH),
        to_signed(4452, D_WIDTH),
        to_signed(4419, D_WIDTH),
        to_signed(4385, D_WIDTH),
        to_signed(4348, D_WIDTH),
        to_signed(4309, D_WIDTH),
        to_signed(4268, D_WIDTH),
        to_signed(4225, D_WIDTH),
        to_signed(4180, D_WIDTH),
        to_signed(4132, D_WIDTH),
        to_signed(4083, D_WIDTH),
        to_signed(4031, D_WIDTH),
        to_signed(3978, D_WIDTH),
        to_signed(3922, D_WIDTH),
        to_signed(3865, D_WIDTH),
        to_signed(3805, D_WIDTH),
        to_signed(3744, D_WIDTH),
        to_signed(3680, D_WIDTH),
        to_signed(3615, D_WIDTH),
        to_signed(3547, D_WIDTH),
        to_signed(3478, D_WIDTH),
        to_signed(3406, D_WIDTH),
        to_signed(3333, D_WIDTH),
        to_signed(3258, D_WIDTH),
        to_signed(3181, D_WIDTH),
        to_signed(3102, D_WIDTH),
        to_signed(3021, D_WIDTH),
        to_signed(2939, D_WIDTH),
        to_signed(2855, D_WIDTH),
        to_signed(2769, D_WIDTH),
        to_signed(2681, D_WIDTH),
        to_signed(2592, D_WIDTH),
        to_signed(2501, D_WIDTH),
        to_signed(2408, D_WIDTH),
        to_signed(2314, D_WIDTH),
        to_signed(2218, D_WIDTH),
        to_signed(2121, D_WIDTH),
        to_signed(2022, D_WIDTH),
        to_signed(1922, D_WIDTH),
        to_signed(1820, D_WIDTH),
        to_signed(1717, D_WIDTH),
        to_signed(1612, D_WIDTH),
        to_signed(1506, D_WIDTH),
        to_signed(1399, D_WIDTH),
        to_signed(1291, D_WIDTH),
        to_signed(1181, D_WIDTH),
        to_signed(1071, D_WIDTH),
        to_signed(959, D_WIDTH),
        to_signed(846, D_WIDTH),
        to_signed(732, D_WIDTH),
        to_signed(617, D_WIDTH),
        to_signed(501, D_WIDTH),
        to_signed(384, D_WIDTH),
        to_signed(266, D_WIDTH),
        to_signed(148, D_WIDTH),
        to_signed(29, D_WIDTH),
        to_signed(-91, D_WIDTH),
        to_signed(-212, D_WIDTH),
        to_signed(-334, D_WIDTH),
        to_signed(-455, D_WIDTH),
        to_signed(-578, D_WIDTH),
        to_signed(-701, D_WIDTH),
        to_signed(-824, D_WIDTH),
        to_signed(-948, D_WIDTH),
        to_signed(-1072, D_WIDTH),
        to_signed(-1197, D_WIDTH),
        to_signed(-1321, D_WIDTH),
        to_signed(-1446, D_WIDTH),
        to_signed(-1571, D_WIDTH),
        to_signed(-1696, D_WIDTH),
        to_signed(-1821, D_WIDTH),
        to_signed(-1946, D_WIDTH),
        to_signed(-2071, D_WIDTH),
        to_signed(-2196, D_WIDTH),
        to_signed(-2320, D_WIDTH),
        to_signed(-2444, D_WIDTH),
        to_signed(-2568, D_WIDTH),
        to_signed(-2692, D_WIDTH),
        to_signed(-2815, D_WIDTH),
        to_signed(-2938, D_WIDTH),
        to_signed(-3060, D_WIDTH),
        to_signed(-3182, D_WIDTH),
        to_signed(-3303, D_WIDTH),
        to_signed(-3423, D_WIDTH),
        to_signed(-3543, D_WIDTH),
        to_signed(-3661, D_WIDTH),
        to_signed(-3779, D_WIDTH),
        to_signed(-3896, D_WIDTH),
        to_signed(-4012, D_WIDTH),
        to_signed(-4127, D_WIDTH),
        to_signed(-4241, D_WIDTH),
        to_signed(-4353, D_WIDTH),
        to_signed(-4465, D_WIDTH),
        to_signed(-4575, D_WIDTH),
        to_signed(-4684, D_WIDTH),
        to_signed(-4791, D_WIDTH),
        to_signed(-4897, D_WIDTH),
        to_signed(-5002, D_WIDTH),
        to_signed(-5105, D_WIDTH),
        to_signed(-5207, D_WIDTH),
        to_signed(-5307, D_WIDTH),
        to_signed(-5405, D_WIDTH),
        to_signed(-5501, D_WIDTH),
        to_signed(-5596, D_WIDTH),
        to_signed(-5689, D_WIDTH),
        to_signed(-5780, D_WIDTH),
        to_signed(-5869, D_WIDTH),
        to_signed(-5955, D_WIDTH),
        to_signed(-6040, D_WIDTH),
        to_signed(-6123, D_WIDTH),
        to_signed(-6204, D_WIDTH),
        to_signed(-6282, D_WIDTH),
        to_signed(-6359, D_WIDTH),
        to_signed(-6433, D_WIDTH),
        to_signed(-6504, D_WIDTH),
        to_signed(-6573, D_WIDTH),
        to_signed(-6640, D_WIDTH),
        to_signed(-6705, D_WIDTH),
        to_signed(-6767, D_WIDTH),
        to_signed(-6826, D_WIDTH),
        to_signed(-6883, D_WIDTH),
        to_signed(-6937, D_WIDTH),
        to_signed(-6988, D_WIDTH),
        to_signed(-7037, D_WIDTH),
        to_signed(-7083, D_WIDTH),
        to_signed(-7126, D_WIDTH),
        to_signed(-7166, D_WIDTH),
        to_signed(-7204, D_WIDTH),
        to_signed(-7239, D_WIDTH),
        to_signed(-7270, D_WIDTH),
        to_signed(-7299, D_WIDTH),
        to_signed(-7325, D_WIDTH),
        to_signed(-7348, D_WIDTH),
        to_signed(-7368, D_WIDTH),
        to_signed(-7384, D_WIDTH),
        to_signed(-7398, D_WIDTH),
        to_signed(-7408, D_WIDTH),
        to_signed(-7416, D_WIDTH),
        to_signed(-7420, D_WIDTH),
        to_signed(-7421, D_WIDTH),
        to_signed(-7419, D_WIDTH),
        to_signed(-7414, D_WIDTH),
        to_signed(-7405, D_WIDTH),
        to_signed(-7393, D_WIDTH),
        to_signed(-7378, D_WIDTH),
        to_signed(-7360, D_WIDTH),
        to_signed(-7338, D_WIDTH),
        to_signed(-7313, D_WIDTH),
        to_signed(-7285, D_WIDTH),
        to_signed(-7253, D_WIDTH),
        to_signed(-7218, D_WIDTH),
        to_signed(-7180, D_WIDTH),
        to_signed(-7138, D_WIDTH),
        to_signed(-7093, D_WIDTH),
        to_signed(-7045, D_WIDTH),
        to_signed(-6993, D_WIDTH),
        to_signed(-6938, D_WIDTH),
        to_signed(-6880, D_WIDTH),
        to_signed(-6818, D_WIDTH),
        to_signed(-6753, D_WIDTH),
        to_signed(-6685, D_WIDTH),
        to_signed(-6614, D_WIDTH),
        to_signed(-6539, D_WIDTH),
        to_signed(-6460, D_WIDTH),
        to_signed(-6379, D_WIDTH),
        to_signed(-6294, D_WIDTH),
        to_signed(-6206, D_WIDTH),
        to_signed(-6115, D_WIDTH),
        to_signed(-6021, D_WIDTH),
        to_signed(-5923, D_WIDTH),
        to_signed(-5823, D_WIDTH),
        to_signed(-5719, D_WIDTH),
        to_signed(-5612, D_WIDTH),
        to_signed(-5502, D_WIDTH),
        to_signed(-5389, D_WIDTH),
        to_signed(-5272, D_WIDTH),
        to_signed(-5153, D_WIDTH),
        to_signed(-5031, D_WIDTH),
        to_signed(-4906, D_WIDTH),
        to_signed(-4778, D_WIDTH),
        to_signed(-4647, D_WIDTH),
        to_signed(-4514, D_WIDTH),
        to_signed(-4377, D_WIDTH),
        to_signed(-4238, D_WIDTH),
        to_signed(-4096, D_WIDTH),
        to_signed(-3952, D_WIDTH),
        to_signed(-3804, D_WIDTH),
        to_signed(-3655, D_WIDTH),
        to_signed(-3503, D_WIDTH),
        to_signed(-3348, D_WIDTH),
        to_signed(-3191, D_WIDTH),
        to_signed(-3031, D_WIDTH),
        to_signed(-2869, D_WIDTH),
        to_signed(-2705, D_WIDTH),
        to_signed(-2539, D_WIDTH),
        to_signed(-2371, D_WIDTH),
        to_signed(-2200, D_WIDTH),
        to_signed(-2028, D_WIDTH),
        to_signed(-1853, D_WIDTH),
        to_signed(-1677, D_WIDTH),
        to_signed(-1499, D_WIDTH),
        to_signed(-1319, D_WIDTH),
        to_signed(-1137, D_WIDTH),
        to_signed(-954, D_WIDTH),
        to_signed(-769, D_WIDTH),
        to_signed(-582, D_WIDTH),
        to_signed(-395, D_WIDTH),
        to_signed(-205, D_WIDTH),
        to_signed(-15, D_WIDTH),
        to_signed(177, D_WIDTH),
        to_signed(370, D_WIDTH),
        to_signed(564, D_WIDTH),
        to_signed(759, D_WIDTH),
        to_signed(955, D_WIDTH),
        to_signed(1151, D_WIDTH),
        to_signed(1349, D_WIDTH),
        to_signed(1547, D_WIDTH),
        to_signed(1746, D_WIDTH),
        to_signed(1945, D_WIDTH),
        to_signed(2145, D_WIDTH),
        to_signed(2345, D_WIDTH),
        to_signed(2545, D_WIDTH),
        to_signed(2746, D_WIDTH),
        to_signed(2946, D_WIDTH),
        to_signed(3147, D_WIDTH),
        to_signed(3348, D_WIDTH),
        to_signed(3548, D_WIDTH),
        to_signed(3748, D_WIDTH),
        to_signed(3948, D_WIDTH),
        to_signed(4148, D_WIDTH),
        to_signed(4347, D_WIDTH),
        to_signed(4545, D_WIDTH),
        to_signed(4743, D_WIDTH),
        to_signed(4940, D_WIDTH),
        to_signed(5136, D_WIDTH),
        to_signed(5331, D_WIDTH),
        to_signed(5526, D_WIDTH),
        to_signed(5719, D_WIDTH),
        to_signed(5911, D_WIDTH),
        to_signed(6101, D_WIDTH),
        to_signed(6290, D_WIDTH),
        to_signed(6478, D_WIDTH),
        to_signed(6664, D_WIDTH),
        to_signed(6849, D_WIDTH),
        to_signed(7031, D_WIDTH),
        to_signed(7212, D_WIDTH),
        to_signed(7391, D_WIDTH),
        to_signed(7568, D_WIDTH),
        to_signed(7743, D_WIDTH),
        to_signed(7916, D_WIDTH),
        to_signed(8086, D_WIDTH),
        to_signed(8255, D_WIDTH),
        to_signed(8420, D_WIDTH),
        to_signed(8583, D_WIDTH),
        to_signed(8744, D_WIDTH),
        to_signed(8902, D_WIDTH),
        to_signed(9057, D_WIDTH),
        to_signed(9209, D_WIDTH),
        to_signed(9358, D_WIDTH),
        to_signed(9504, D_WIDTH),
        to_signed(9647, D_WIDTH),
        to_signed(9787, D_WIDTH),
        to_signed(9923, D_WIDTH),
        to_signed(10056, D_WIDTH),
        to_signed(10186, D_WIDTH),
        to_signed(10312, D_WIDTH),
        to_signed(10435, D_WIDTH),
        to_signed(10554, D_WIDTH),
        to_signed(10669, D_WIDTH),
        to_signed(10780, D_WIDTH),
        to_signed(10888, D_WIDTH),
        to_signed(10991, D_WIDTH),
        to_signed(11091, D_WIDTH),
        to_signed(11186, D_WIDTH),
        to_signed(11277, D_WIDTH),
        to_signed(11364, D_WIDTH),
        to_signed(11447, D_WIDTH),
        to_signed(11525, D_WIDTH),
        to_signed(11599, D_WIDTH),
        to_signed(11668, D_WIDTH),
        to_signed(11733, D_WIDTH),
        to_signed(11793, D_WIDTH),
        to_signed(11848, D_WIDTH),
        to_signed(11899, D_WIDTH),
        to_signed(11945, D_WIDTH),
        to_signed(11986, D_WIDTH),
        to_signed(12022, D_WIDTH),
        to_signed(12054, D_WIDTH),
        to_signed(12080, D_WIDTH),
        to_signed(12101, D_WIDTH),
        to_signed(12117, D_WIDTH),
        to_signed(12128, D_WIDTH),
        to_signed(12134, D_WIDTH),
        to_signed(12135, D_WIDTH),
        to_signed(12131, D_WIDTH),
        to_signed(12121, D_WIDTH),
        to_signed(12106, D_WIDTH),
        to_signed(12085, D_WIDTH),
        to_signed(12060, D_WIDTH),
        to_signed(12029, D_WIDTH),
        to_signed(11992, D_WIDTH),
        to_signed(11950, D_WIDTH),
        to_signed(11903, D_WIDTH),
        to_signed(11850, D_WIDTH),
        to_signed(11792, D_WIDTH),
        to_signed(11728, D_WIDTH),
        to_signed(11658, D_WIDTH),
        to_signed(11583, D_WIDTH),
        to_signed(11503, D_WIDTH),
        to_signed(11417, D_WIDTH),
        to_signed(11326, D_WIDTH),
        to_signed(11229, D_WIDTH),
        to_signed(11126, D_WIDTH),
        to_signed(11018, D_WIDTH),
        to_signed(10904, D_WIDTH),
        to_signed(10785, D_WIDTH),
        to_signed(10660, D_WIDTH),
        to_signed(10530, D_WIDTH),
        to_signed(10395, D_WIDTH),
        to_signed(10254, D_WIDTH),
        to_signed(10107, D_WIDTH),
        to_signed(9955, D_WIDTH),
        to_signed(9798, D_WIDTH),
        to_signed(9635, D_WIDTH),
        to_signed(9467, D_WIDTH),
        to_signed(9293, D_WIDTH),
        to_signed(9115, D_WIDTH),
        to_signed(8931, D_WIDTH),
        to_signed(8741, D_WIDTH),
        to_signed(8547, D_WIDTH),
        to_signed(8348, D_WIDTH),
        to_signed(8143, D_WIDTH),
        to_signed(7934, D_WIDTH),
        to_signed(7719, D_WIDTH),
        to_signed(7499, D_WIDTH),
        to_signed(7275, D_WIDTH),
        to_signed(7046, D_WIDTH),
        to_signed(6812, D_WIDTH),
        to_signed(6573, D_WIDTH),
        to_signed(6330, D_WIDTH),
        to_signed(6082, D_WIDTH),
        to_signed(5830, D_WIDTH),
        to_signed(5573, D_WIDTH),
        to_signed(5312, D_WIDTH),
        to_signed(5047, D_WIDTH),
        to_signed(4777, D_WIDTH),
        to_signed(4504, D_WIDTH),
        to_signed(4226, D_WIDTH),
        to_signed(3944, D_WIDTH),
        to_signed(3659, D_WIDTH),
        to_signed(3370, D_WIDTH),
        to_signed(3077, D_WIDTH),
        to_signed(2780, D_WIDTH),
        to_signed(2480, D_WIDTH),
        to_signed(2177, D_WIDTH),
        to_signed(1870, D_WIDTH),
        to_signed(1560, D_WIDTH),
        to_signed(1247, D_WIDTH),
        to_signed(931, D_WIDTH),
        to_signed(612, D_WIDTH),
        to_signed(290, D_WIDTH),
        to_signed(-34, D_WIDTH),
        to_signed(-361, D_WIDTH),
        to_signed(-690, D_WIDTH),
        to_signed(-1022, D_WIDTH),
        to_signed(-1355, D_WIDTH),
        to_signed(-1691, D_WIDTH),
        to_signed(-2029, D_WIDTH),
        to_signed(-2369, D_WIDTH),
        to_signed(-2710, D_WIDTH),
        to_signed(-3053, D_WIDTH),
        to_signed(-3397, D_WIDTH),
        to_signed(-3743, D_WIDTH),
        to_signed(-4090, D_WIDTH),
        to_signed(-4437, D_WIDTH),
        to_signed(-4786, D_WIDTH),
        to_signed(-5136, D_WIDTH),
        to_signed(-5486, D_WIDTH),
        to_signed(-5837, D_WIDTH),
        to_signed(-6188, D_WIDTH),
        to_signed(-6539, D_WIDTH),
        to_signed(-6890, D_WIDTH),
        to_signed(-7242, D_WIDTH),
        to_signed(-7593, D_WIDTH),
        to_signed(-7943, D_WIDTH),
        to_signed(-8293, D_WIDTH),
        to_signed(-8643, D_WIDTH),
        to_signed(-8992, D_WIDTH),
        to_signed(-9339, D_WIDTH),
        to_signed(-9686, D_WIDTH),
        to_signed(-10032, D_WIDTH),
        to_signed(-10375, D_WIDTH),
        to_signed(-10718, D_WIDTH),
        to_signed(-11059, D_WIDTH),
        to_signed(-11397, D_WIDTH),
        to_signed(-11734, D_WIDTH),
        to_signed(-12069, D_WIDTH),
        to_signed(-12401, D_WIDTH),
        to_signed(-12731, D_WIDTH),
        to_signed(-13058, D_WIDTH),
        to_signed(-13383, D_WIDTH),
        to_signed(-13704, D_WIDTH),
        to_signed(-14022, D_WIDTH),
        to_signed(-14338, D_WIDTH),
        to_signed(-14649, D_WIDTH),
        to_signed(-14957, D_WIDTH),
        to_signed(-15261, D_WIDTH),
        to_signed(-15562, D_WIDTH),
        to_signed(-15858, D_WIDTH),
        to_signed(-16150, D_WIDTH),
        to_signed(-16438, D_WIDTH),
        to_signed(-16721, D_WIDTH),
        to_signed(-17000, D_WIDTH),
        to_signed(-17274, D_WIDTH),
        to_signed(-17543, D_WIDTH),
        to_signed(-17806, D_WIDTH),
        to_signed(-18064, D_WIDTH),
        to_signed(-18317, D_WIDTH),
        to_signed(-18565, D_WIDTH),
        to_signed(-18806, D_WIDTH),
        to_signed(-19042, D_WIDTH),
        to_signed(-19272, D_WIDTH),
        to_signed(-19495, D_WIDTH),
        to_signed(-19712, D_WIDTH),
        to_signed(-19923, D_WIDTH),
        to_signed(-20127, D_WIDTH),
        to_signed(-20324, D_WIDTH),
        to_signed(-20514, D_WIDTH),
        to_signed(-20697, D_WIDTH),
        to_signed(-20873, D_WIDTH),
        to_signed(-21042, D_WIDTH),
        to_signed(-21203, D_WIDTH),
        to_signed(-21357, D_WIDTH),
        to_signed(-21503, D_WIDTH),
        to_signed(-21641, D_WIDTH),
        to_signed(-21771, D_WIDTH),
        to_signed(-21893, D_WIDTH),
        to_signed(-22006, D_WIDTH),
        to_signed(-22111, D_WIDTH),
        to_signed(-22208, D_WIDTH),
        to_signed(-22296, D_WIDTH),
        to_signed(-22375, D_WIDTH),
        to_signed(-22446, D_WIDTH),
        to_signed(-22507, D_WIDTH),
        to_signed(-22560, D_WIDTH),
        to_signed(-22603, D_WIDTH),
        to_signed(-22637, D_WIDTH),
        to_signed(-22661, D_WIDTH),
        to_signed(-22676, D_WIDTH),
        to_signed(-22681, D_WIDTH),
        to_signed(-22677, D_WIDTH),
        to_signed(-22662, D_WIDTH),
        to_signed(-22638, D_WIDTH),
        to_signed(-22604, D_WIDTH),
        to_signed(-22559, D_WIDTH),
        to_signed(-22505, D_WIDTH),
        to_signed(-22440, D_WIDTH),
        to_signed(-22365, D_WIDTH),
        to_signed(-22279, D_WIDTH),
        to_signed(-22183, D_WIDTH),
        to_signed(-22076, D_WIDTH),
        to_signed(-21959, D_WIDTH),
        to_signed(-21830, D_WIDTH),
        to_signed(-21691, D_WIDTH),
        to_signed(-21542, D_WIDTH),
        to_signed(-21381, D_WIDTH),
        to_signed(-21209, D_WIDTH),
        to_signed(-21027, D_WIDTH),
        to_signed(-20833, D_WIDTH),
        to_signed(-20628, D_WIDTH),
        to_signed(-20412, D_WIDTH),
        to_signed(-20185, D_WIDTH),
        to_signed(-19946, D_WIDTH),
        to_signed(-19696, D_WIDTH),
        to_signed(-19435, D_WIDTH),
        to_signed(-19163, D_WIDTH),
        to_signed(-18879, D_WIDTH),
        to_signed(-18584, D_WIDTH),
        to_signed(-18277, D_WIDTH),
        to_signed(-17959, D_WIDTH),
        to_signed(-17630, D_WIDTH),
        to_signed(-17289, D_WIDTH),
        to_signed(-16937, D_WIDTH),
        to_signed(-16573, D_WIDTH),
        to_signed(-16198, D_WIDTH),
        to_signed(-15812, D_WIDTH),
        to_signed(-15414, D_WIDTH),
        to_signed(-15004, D_WIDTH),
        to_signed(-14584, D_WIDTH),
        to_signed(-14152, D_WIDTH),
        to_signed(-13708, D_WIDTH),
        to_signed(-13253, D_WIDTH),
        to_signed(-12787, D_WIDTH),
        to_signed(-12310, D_WIDTH),
        to_signed(-11822, D_WIDTH),
        to_signed(-11322, D_WIDTH),
        to_signed(-10812, D_WIDTH),
        to_signed(-10290, D_WIDTH),
        to_signed(-9757, D_WIDTH),
        to_signed(-9213, D_WIDTH),
        to_signed(-8659, D_WIDTH),
        to_signed(-8093, D_WIDTH),
        to_signed(-7517, D_WIDTH),
        to_signed(-6930, D_WIDTH),
        to_signed(-6332, D_WIDTH),
        to_signed(-5724, D_WIDTH),
        to_signed(-5105, D_WIDTH),
        to_signed(-4476, D_WIDTH),
        to_signed(-3837, D_WIDTH),
        to_signed(-3187, D_WIDTH),
        to_signed(-2528, D_WIDTH),
        to_signed(-1858, D_WIDTH),
        to_signed(-1179, D_WIDTH),
        to_signed(-489, D_WIDTH),
        to_signed(210, D_WIDTH),
        to_signed(919, D_WIDTH),
        to_signed(1637, D_WIDTH),
        to_signed(2364, D_WIDTH),
        to_signed(3101, D_WIDTH),
        to_signed(3847, D_WIDTH),
        to_signed(4602, D_WIDTH),
        to_signed(5366, D_WIDTH),
        to_signed(6138, D_WIDTH),
        to_signed(6919, D_WIDTH),
        to_signed(7709, D_WIDTH),
        to_signed(8507, D_WIDTH),
        to_signed(9313, D_WIDTH),
        to_signed(10127, D_WIDTH),
        to_signed(10949, D_WIDTH),
        to_signed(11779, D_WIDTH),
        to_signed(12616, D_WIDTH),
        to_signed(13460, D_WIDTH),
        to_signed(14312, D_WIDTH),
        to_signed(15171, D_WIDTH),
        to_signed(16037, D_WIDTH),
        to_signed(16909, D_WIDTH),
        to_signed(17788, D_WIDTH),
        to_signed(18674, D_WIDTH),
        to_signed(19565, D_WIDTH),
        to_signed(20463, D_WIDTH),
        to_signed(21366, D_WIDTH),
        to_signed(22275, D_WIDTH),
        to_signed(23190, D_WIDTH),
        to_signed(24110, D_WIDTH),
        to_signed(25035, D_WIDTH),
        to_signed(25964, D_WIDTH),
        to_signed(26899, D_WIDTH),
        to_signed(27838, D_WIDTH),
        to_signed(28781, D_WIDTH),
        to_signed(29728, D_WIDTH),
        to_signed(30679, D_WIDTH),
        to_signed(31634, D_WIDTH),
        to_signed(32593, D_WIDTH),
        to_signed(33554, D_WIDTH),
        to_signed(34519, D_WIDTH),
        to_signed(35486, D_WIDTH),
        to_signed(36456, D_WIDTH),
        to_signed(37428, D_WIDTH),
        to_signed(38403, D_WIDTH),
        to_signed(39380, D_WIDTH),
        to_signed(40358, D_WIDTH),
        to_signed(41337, D_WIDTH),
        to_signed(42318, D_WIDTH),
        to_signed(43301, D_WIDTH),
        to_signed(44283, D_WIDTH),
        to_signed(45267, D_WIDTH),
        to_signed(46251, D_WIDTH),
        to_signed(47235, D_WIDTH),
        to_signed(48219, D_WIDTH),
        to_signed(49203, D_WIDTH),
        to_signed(50186, D_WIDTH),
        to_signed(51168, D_WIDTH),
        to_signed(52150, D_WIDTH),
        to_signed(53130, D_WIDTH),
        to_signed(54108, D_WIDTH),
        to_signed(55085, D_WIDTH),
        to_signed(56061, D_WIDTH),
        to_signed(57033, D_WIDTH),
        to_signed(58004, D_WIDTH),
        to_signed(58972, D_WIDTH),
        to_signed(59937, D_WIDTH),
        to_signed(60899, D_WIDTH),
        to_signed(61858, D_WIDTH),
        to_signed(62813, D_WIDTH),
        to_signed(63764, D_WIDTH),
        to_signed(64711, D_WIDTH),
        to_signed(65654, D_WIDTH),
        to_signed(66593, D_WIDTH),
        to_signed(67527, D_WIDTH),
        to_signed(68456, D_WIDTH),
        to_signed(69379, D_WIDTH),
        to_signed(70298, D_WIDTH),
        to_signed(71211, D_WIDTH),
        to_signed(72117, D_WIDTH),
        to_signed(73018, D_WIDTH),
        to_signed(73913, D_WIDTH),
        to_signed(74801, D_WIDTH),
        to_signed(75682, D_WIDTH),
        to_signed(76557, D_WIDTH),
        to_signed(77424, D_WIDTH),
        to_signed(78283, D_WIDTH),
        to_signed(79136, D_WIDTH),
        to_signed(79980, D_WIDTH),
        to_signed(80816, D_WIDTH),
        to_signed(81644, D_WIDTH),
        to_signed(82464, D_WIDTH),
        to_signed(83275, D_WIDTH),
        to_signed(84077, D_WIDTH),
        to_signed(84870, D_WIDTH),
        to_signed(85654, D_WIDTH),
        to_signed(86428, D_WIDTH),
        to_signed(87193, D_WIDTH),
        to_signed(87948, D_WIDTH),
        to_signed(88692, D_WIDTH),
        to_signed(89427, D_WIDTH),
        to_signed(90151, D_WIDTH),
        to_signed(90865, D_WIDTH),
        to_signed(91567, D_WIDTH),
        to_signed(92259, D_WIDTH),
        to_signed(92940, D_WIDTH),
        to_signed(93609, D_WIDTH),
        to_signed(94266, D_WIDTH),
        to_signed(94913, D_WIDTH),
        to_signed(95547, D_WIDTH),
        to_signed(96169, D_WIDTH),
        to_signed(96779, D_WIDTH),
        to_signed(97377, D_WIDTH),
        to_signed(97962, D_WIDTH),
        to_signed(98535, D_WIDTH),
        to_signed(99095, D_WIDTH),
        to_signed(99642, D_WIDTH),
        to_signed(100176, D_WIDTH),
        to_signed(100697, D_WIDTH),
        to_signed(101204, D_WIDTH),
        to_signed(101698, D_WIDTH),
        to_signed(102178, D_WIDTH),
        to_signed(102645, D_WIDTH),
        to_signed(103098, D_WIDTH),
        to_signed(103537, D_WIDTH),
        to_signed(103962, D_WIDTH),
        to_signed(104372, D_WIDTH),
        to_signed(104769, D_WIDTH),
        to_signed(105151, D_WIDTH),
        to_signed(105518, D_WIDTH),
        to_signed(105871, D_WIDTH),
        to_signed(106209, D_WIDTH),
        to_signed(106533, D_WIDTH),
        to_signed(106841, D_WIDTH),
        to_signed(107135, D_WIDTH),
        to_signed(107414, D_WIDTH),
        to_signed(107677, D_WIDTH),
        to_signed(107926, D_WIDTH),
        to_signed(108159, D_WIDTH),
        to_signed(108377, D_WIDTH),
        to_signed(108580, D_WIDTH),
        to_signed(108767, D_WIDTH),
        to_signed(108939, D_WIDTH),
        to_signed(109095, D_WIDTH),
        to_signed(109236, D_WIDTH),
        to_signed(109361, D_WIDTH),
        to_signed(109471, D_WIDTH),
        to_signed(109565, D_WIDTH),
        to_signed(109643, D_WIDTH),
        to_signed(109706, D_WIDTH),
        to_signed(109753, D_WIDTH),
        to_signed(109785, D_WIDTH),
        to_signed(109800, D_WIDTH),

        -- 2048 - 1920 = 128 padding works
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH)
    );

begin

    process(clk)
    begin
        if rising_edge(clk) then
            if clk_en = '1' then
                data <= coeff_list(to_integer(addr));
            end if;
        end if;
    end process;

end rtl;
