library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity coeff_rom is
    generic(
        A_WIDTH : integer;
        D_WIDTH : integer
        );
    port (
        clk    : in  std_logic;
        clk_en : in  std_logic;
        addr   : in  unsigned(A_WIDTH - 1 downto 0);
        data   : out signed(D_WIDTH - 1 downto 0)
        );
end;

architecture rtl of coeff_rom is

    type t_coeff_list is array(0 to 2 ** A_WIDTH - 1) of
        signed(D_WIDTH - 1 downto 0);

    signal coeff_list : t_coeff_list := (
        to_signed(-108, D_WIDTH),
        to_signed(-107, D_WIDTH),
        to_signed(-105, D_WIDTH),
        to_signed(-104, D_WIDTH),
        to_signed(-102, D_WIDTH),
        to_signed(-100, D_WIDTH),
        to_signed(-99, D_WIDTH),
        to_signed(-97, D_WIDTH),
        to_signed(-95, D_WIDTH),
        to_signed(-94, D_WIDTH),
        to_signed(-92, D_WIDTH),
        to_signed(-90, D_WIDTH),
        to_signed(-88, D_WIDTH),
        to_signed(-86, D_WIDTH),
        to_signed(-84, D_WIDTH),
        to_signed(-82, D_WIDTH),
        to_signed(-80, D_WIDTH),
        to_signed(-78, D_WIDTH),
        to_signed(-76, D_WIDTH),
        to_signed(-74, D_WIDTH),
        to_signed(-72, D_WIDTH),
        to_signed(-70, D_WIDTH),
        to_signed(-68, D_WIDTH),
        to_signed(-65, D_WIDTH),
        to_signed(-63, D_WIDTH),
        to_signed(-61, D_WIDTH),
        to_signed(-59, D_WIDTH),
        to_signed(-56, D_WIDTH),
        to_signed(-54, D_WIDTH),
        to_signed(-52, D_WIDTH),
        to_signed(-49, D_WIDTH),
        to_signed(-47, D_WIDTH),
        to_signed(-45, D_WIDTH),
        to_signed(-42, D_WIDTH),
        to_signed(-40, D_WIDTH),
        to_signed(-37, D_WIDTH),
        to_signed(-35, D_WIDTH),
        to_signed(-32, D_WIDTH),
        to_signed(-30, D_WIDTH),
        to_signed(-27, D_WIDTH),
        to_signed(-25, D_WIDTH),
        to_signed(-22, D_WIDTH),
        to_signed(-19, D_WIDTH),
        to_signed(-17, D_WIDTH),
        to_signed(-14, D_WIDTH),
        to_signed(-12, D_WIDTH),
        to_signed(-9, D_WIDTH),
        to_signed(-6, D_WIDTH),
        to_signed(-4, D_WIDTH),
        to_signed(-1, D_WIDTH),
        to_signed(2, D_WIDTH),
        to_signed(4, D_WIDTH),
        to_signed(7, D_WIDTH),
        to_signed(10, D_WIDTH),
        to_signed(13, D_WIDTH),
        to_signed(15, D_WIDTH),
        to_signed(18, D_WIDTH),
        to_signed(21, D_WIDTH),
        to_signed(23, D_WIDTH),
        to_signed(26, D_WIDTH),
        to_signed(29, D_WIDTH),
        to_signed(32, D_WIDTH),
        to_signed(34, D_WIDTH),
        to_signed(37, D_WIDTH),
        to_signed(40, D_WIDTH),
        to_signed(42, D_WIDTH),
        to_signed(45, D_WIDTH),
        to_signed(48, D_WIDTH),
        to_signed(51, D_WIDTH),
        to_signed(53, D_WIDTH),
        to_signed(56, D_WIDTH),
        to_signed(59, D_WIDTH),
        to_signed(61, D_WIDTH),
        to_signed(64, D_WIDTH),
        to_signed(67, D_WIDTH),
        to_signed(69, D_WIDTH),
        to_signed(72, D_WIDTH),
        to_signed(74, D_WIDTH),
        to_signed(77, D_WIDTH),
        to_signed(79, D_WIDTH),
        to_signed(82, D_WIDTH),
        to_signed(85, D_WIDTH),
        to_signed(87, D_WIDTH),
        to_signed(90, D_WIDTH),
        to_signed(92, D_WIDTH),
        to_signed(94, D_WIDTH),
        to_signed(97, D_WIDTH),
        to_signed(99, D_WIDTH),
        to_signed(102, D_WIDTH),
        to_signed(104, D_WIDTH),
        to_signed(106, D_WIDTH),
        to_signed(109, D_WIDTH),
        to_signed(111, D_WIDTH),
        to_signed(113, D_WIDTH),
        to_signed(115, D_WIDTH),
        to_signed(118, D_WIDTH),
        to_signed(120, D_WIDTH),
        to_signed(122, D_WIDTH),
        to_signed(124, D_WIDTH),
        to_signed(126, D_WIDTH),
        to_signed(128, D_WIDTH),
        to_signed(130, D_WIDTH),
        to_signed(132, D_WIDTH),
        to_signed(134, D_WIDTH),
        to_signed(136, D_WIDTH),
        to_signed(138, D_WIDTH),
        to_signed(140, D_WIDTH),
        to_signed(141, D_WIDTH),
        to_signed(143, D_WIDTH),
        to_signed(145, D_WIDTH),
        to_signed(147, D_WIDTH),
        to_signed(148, D_WIDTH),
        to_signed(150, D_WIDTH),
        to_signed(151, D_WIDTH),
        to_signed(153, D_WIDTH),
        to_signed(154, D_WIDTH),
        to_signed(156, D_WIDTH),
        to_signed(157, D_WIDTH),
        to_signed(158, D_WIDTH),
        to_signed(160, D_WIDTH),
        to_signed(161, D_WIDTH),
        to_signed(162, D_WIDTH),
        to_signed(163, D_WIDTH),
        to_signed(164, D_WIDTH),
        to_signed(165, D_WIDTH),
        to_signed(166, D_WIDTH),
        to_signed(167, D_WIDTH),
        to_signed(168, D_WIDTH),
        to_signed(169, D_WIDTH),
        to_signed(169, D_WIDTH),
        to_signed(170, D_WIDTH),
        to_signed(171, D_WIDTH),
        to_signed(171, D_WIDTH),
        to_signed(172, D_WIDTH),
        to_signed(172, D_WIDTH),
        to_signed(173, D_WIDTH),
        to_signed(173, D_WIDTH),
        to_signed(174, D_WIDTH),
        to_signed(174, D_WIDTH),
        to_signed(174, D_WIDTH),
        to_signed(174, D_WIDTH),
        to_signed(174, D_WIDTH),
        to_signed(174, D_WIDTH),
        to_signed(174, D_WIDTH),
        to_signed(174, D_WIDTH),
        to_signed(174, D_WIDTH),
        to_signed(174, D_WIDTH),
        to_signed(173, D_WIDTH),
        to_signed(173, D_WIDTH),
        to_signed(173, D_WIDTH),
        to_signed(172, D_WIDTH),
        to_signed(172, D_WIDTH),
        to_signed(171, D_WIDTH),
        to_signed(171, D_WIDTH),
        to_signed(170, D_WIDTH),
        to_signed(169, D_WIDTH),
        to_signed(168, D_WIDTH),
        to_signed(167, D_WIDTH),
        to_signed(166, D_WIDTH),
        to_signed(165, D_WIDTH),
        to_signed(164, D_WIDTH),
        to_signed(163, D_WIDTH),
        to_signed(162, D_WIDTH),
        to_signed(161, D_WIDTH),
        to_signed(159, D_WIDTH),
        to_signed(158, D_WIDTH),
        to_signed(156, D_WIDTH),
        to_signed(155, D_WIDTH),
        to_signed(153, D_WIDTH),
        to_signed(152, D_WIDTH),
        to_signed(150, D_WIDTH),
        to_signed(148, D_WIDTH),
        to_signed(146, D_WIDTH),
        to_signed(145, D_WIDTH),
        to_signed(143, D_WIDTH),
        to_signed(141, D_WIDTH),
        to_signed(139, D_WIDTH),
        to_signed(136, D_WIDTH),
        to_signed(134, D_WIDTH),
        to_signed(132, D_WIDTH),
        to_signed(130, D_WIDTH),
        to_signed(127, D_WIDTH),
        to_signed(125, D_WIDTH),
        to_signed(122, D_WIDTH),
        to_signed(120, D_WIDTH),
        to_signed(117, D_WIDTH),
        to_signed(115, D_WIDTH),
        to_signed(112, D_WIDTH),
        to_signed(109, D_WIDTH),
        to_signed(106, D_WIDTH),
        to_signed(104, D_WIDTH),
        to_signed(101, D_WIDTH),
        to_signed(98, D_WIDTH),
        to_signed(95, D_WIDTH),
        to_signed(92, D_WIDTH),
        to_signed(88, D_WIDTH),
        to_signed(85, D_WIDTH),
        to_signed(82, D_WIDTH),
        to_signed(79, D_WIDTH),
        to_signed(75, D_WIDTH),
        to_signed(72, D_WIDTH),
        to_signed(69, D_WIDTH),
        to_signed(65, D_WIDTH),
        to_signed(62, D_WIDTH),
        to_signed(58, D_WIDTH),
        to_signed(55, D_WIDTH),
        to_signed(51, D_WIDTH),
        to_signed(47, D_WIDTH),
        to_signed(44, D_WIDTH),
        to_signed(40, D_WIDTH),
        to_signed(36, D_WIDTH),
        to_signed(32, D_WIDTH),
        to_signed(28, D_WIDTH),
        to_signed(24, D_WIDTH),
        to_signed(21, D_WIDTH),
        to_signed(17, D_WIDTH),
        to_signed(13, D_WIDTH),
        to_signed(9, D_WIDTH),
        to_signed(5, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(-4, D_WIDTH),
        to_signed(-8, D_WIDTH),
        to_signed(-12, D_WIDTH),
        to_signed(-16, D_WIDTH),
        to_signed(-20, D_WIDTH),
        to_signed(-25, D_WIDTH),
        to_signed(-29, D_WIDTH),
        to_signed(-33, D_WIDTH),
        to_signed(-37, D_WIDTH),
        to_signed(-42, D_WIDTH),
        to_signed(-46, D_WIDTH),
        to_signed(-50, D_WIDTH),
        to_signed(-54, D_WIDTH),
        to_signed(-59, D_WIDTH),
        to_signed(-63, D_WIDTH),
        to_signed(-67, D_WIDTH),
        to_signed(-72, D_WIDTH),
        to_signed(-76, D_WIDTH),
        to_signed(-80, D_WIDTH),
        to_signed(-85, D_WIDTH),
        to_signed(-89, D_WIDTH),
        to_signed(-94, D_WIDTH),
        to_signed(-98, D_WIDTH),
        to_signed(-102, D_WIDTH),
        to_signed(-107, D_WIDTH),
        to_signed(-111, D_WIDTH),
        to_signed(-115, D_WIDTH),
        to_signed(-119, D_WIDTH),
        to_signed(-124, D_WIDTH),
        to_signed(-128, D_WIDTH),
        to_signed(-132, D_WIDTH),
        to_signed(-137, D_WIDTH),
        to_signed(-141, D_WIDTH),
        to_signed(-145, D_WIDTH),
        to_signed(-149, D_WIDTH),
        to_signed(-153, D_WIDTH),
        to_signed(-157, D_WIDTH),
        to_signed(-161, D_WIDTH),
        to_signed(-166, D_WIDTH),
        to_signed(-170, D_WIDTH),
        to_signed(-174, D_WIDTH),
        to_signed(-178, D_WIDTH),
        to_signed(-182, D_WIDTH),
        to_signed(-185, D_WIDTH),
        to_signed(-189, D_WIDTH),
        to_signed(-193, D_WIDTH),
        to_signed(-197, D_WIDTH),
        to_signed(-201, D_WIDTH),
        to_signed(-204, D_WIDTH),
        to_signed(-208, D_WIDTH),
        to_signed(-211, D_WIDTH),
        to_signed(-215, D_WIDTH),
        to_signed(-219, D_WIDTH),
        to_signed(-222, D_WIDTH),
        to_signed(-225, D_WIDTH),
        to_signed(-229, D_WIDTH),
        to_signed(-232, D_WIDTH),
        to_signed(-235, D_WIDTH),
        to_signed(-238, D_WIDTH),
        to_signed(-241, D_WIDTH),
        to_signed(-244, D_WIDTH),
        to_signed(-247, D_WIDTH),
        to_signed(-250, D_WIDTH),
        to_signed(-253, D_WIDTH),
        to_signed(-256, D_WIDTH),
        to_signed(-258, D_WIDTH),
        to_signed(-261, D_WIDTH),
        to_signed(-264, D_WIDTH),
        to_signed(-266, D_WIDTH),
        to_signed(-268, D_WIDTH),
        to_signed(-271, D_WIDTH),
        to_signed(-273, D_WIDTH),
        to_signed(-275, D_WIDTH),
        to_signed(-277, D_WIDTH),
        to_signed(-279, D_WIDTH),
        to_signed(-281, D_WIDTH),
        to_signed(-283, D_WIDTH),
        to_signed(-284, D_WIDTH),
        to_signed(-286, D_WIDTH),
        to_signed(-288, D_WIDTH),
        to_signed(-289, D_WIDTH),
        to_signed(-290, D_WIDTH),
        to_signed(-292, D_WIDTH),
        to_signed(-293, D_WIDTH),
        to_signed(-294, D_WIDTH),
        to_signed(-295, D_WIDTH),
        to_signed(-296, D_WIDTH),
        to_signed(-297, D_WIDTH),
        to_signed(-297, D_WIDTH),
        to_signed(-298, D_WIDTH),
        to_signed(-298, D_WIDTH),
        to_signed(-299, D_WIDTH),
        to_signed(-299, D_WIDTH),
        to_signed(-299, D_WIDTH),
        to_signed(-299, D_WIDTH),
        to_signed(-299, D_WIDTH),
        to_signed(-299, D_WIDTH),
        to_signed(-299, D_WIDTH),
        to_signed(-298, D_WIDTH),
        to_signed(-298, D_WIDTH),
        to_signed(-297, D_WIDTH),
        to_signed(-296, D_WIDTH),
        to_signed(-296, D_WIDTH),
        to_signed(-295, D_WIDTH),
        to_signed(-294, D_WIDTH),
        to_signed(-293, D_WIDTH),
        to_signed(-291, D_WIDTH),
        to_signed(-290, D_WIDTH),
        to_signed(-288, D_WIDTH),
        to_signed(-287, D_WIDTH),
        to_signed(-285, D_WIDTH),
        to_signed(-283, D_WIDTH),
        to_signed(-281, D_WIDTH),
        to_signed(-279, D_WIDTH),
        to_signed(-277, D_WIDTH),
        to_signed(-275, D_WIDTH),
        to_signed(-273, D_WIDTH),
        to_signed(-270, D_WIDTH),
        to_signed(-268, D_WIDTH),
        to_signed(-265, D_WIDTH),
        to_signed(-262, D_WIDTH),
        to_signed(-259, D_WIDTH),
        to_signed(-256, D_WIDTH),
        to_signed(-253, D_WIDTH),
        to_signed(-249, D_WIDTH),
        to_signed(-246, D_WIDTH),
        to_signed(-243, D_WIDTH),
        to_signed(-239, D_WIDTH),
        to_signed(-235, D_WIDTH),
        to_signed(-231, D_WIDTH),
        to_signed(-227, D_WIDTH),
        to_signed(-223, D_WIDTH),
        to_signed(-219, D_WIDTH),
        to_signed(-215, D_WIDTH),
        to_signed(-211, D_WIDTH),
        to_signed(-206, D_WIDTH),
        to_signed(-202, D_WIDTH),
        to_signed(-197, D_WIDTH),
        to_signed(-192, D_WIDTH),
        to_signed(-187, D_WIDTH),
        to_signed(-182, D_WIDTH),
        to_signed(-177, D_WIDTH),
        to_signed(-172, D_WIDTH),
        to_signed(-167, D_WIDTH),
        to_signed(-161, D_WIDTH),
        to_signed(-156, D_WIDTH),
        to_signed(-150, D_WIDTH),
        to_signed(-145, D_WIDTH),
        to_signed(-139, D_WIDTH),
        to_signed(-133, D_WIDTH),
        to_signed(-127, D_WIDTH),
        to_signed(-121, D_WIDTH),
        to_signed(-115, D_WIDTH),
        to_signed(-109, D_WIDTH),
        to_signed(-102, D_WIDTH),
        to_signed(-96, D_WIDTH),
        to_signed(-90, D_WIDTH),
        to_signed(-83, D_WIDTH),
        to_signed(-77, D_WIDTH),
        to_signed(-70, D_WIDTH),
        to_signed(-63, D_WIDTH),
        to_signed(-56, D_WIDTH),
        to_signed(-50, D_WIDTH),
        to_signed(-43, D_WIDTH),
        to_signed(-36, D_WIDTH),
        to_signed(-29, D_WIDTH),
        to_signed(-21, D_WIDTH),
        to_signed(-14, D_WIDTH),
        to_signed(-7, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(8, D_WIDTH),
        to_signed(15, D_WIDTH),
        to_signed(22, D_WIDTH),
        to_signed(30, D_WIDTH),
        to_signed(37, D_WIDTH),
        to_signed(45, D_WIDTH),
        to_signed(52, D_WIDTH),
        to_signed(60, D_WIDTH),
        to_signed(68, D_WIDTH),
        to_signed(75, D_WIDTH),
        to_signed(83, D_WIDTH),
        to_signed(91, D_WIDTH),
        to_signed(98, D_WIDTH),
        to_signed(106, D_WIDTH),
        to_signed(114, D_WIDTH),
        to_signed(122, D_WIDTH),
        to_signed(130, D_WIDTH),
        to_signed(137, D_WIDTH),
        to_signed(145, D_WIDTH),
        to_signed(153, D_WIDTH),
        to_signed(161, D_WIDTH),
        to_signed(169, D_WIDTH),
        to_signed(176, D_WIDTH),
        to_signed(184, D_WIDTH),
        to_signed(192, D_WIDTH),
        to_signed(200, D_WIDTH),
        to_signed(207, D_WIDTH),
        to_signed(215, D_WIDTH),
        to_signed(223, D_WIDTH),
        to_signed(231, D_WIDTH),
        to_signed(238, D_WIDTH),
        to_signed(246, D_WIDTH),
        to_signed(253, D_WIDTH),
        to_signed(261, D_WIDTH),
        to_signed(268, D_WIDTH),
        to_signed(276, D_WIDTH),
        to_signed(283, D_WIDTH),
        to_signed(291, D_WIDTH),
        to_signed(298, D_WIDTH),
        to_signed(305, D_WIDTH),
        to_signed(312, D_WIDTH),
        to_signed(320, D_WIDTH),
        to_signed(327, D_WIDTH),
        to_signed(334, D_WIDTH),
        to_signed(341, D_WIDTH),
        to_signed(347, D_WIDTH),
        to_signed(354, D_WIDTH),
        to_signed(361, D_WIDTH),
        to_signed(368, D_WIDTH),
        to_signed(374, D_WIDTH),
        to_signed(380, D_WIDTH),
        to_signed(387, D_WIDTH),
        to_signed(393, D_WIDTH),
        to_signed(399, D_WIDTH),
        to_signed(405, D_WIDTH),
        to_signed(411, D_WIDTH),
        to_signed(417, D_WIDTH),
        to_signed(423, D_WIDTH),
        to_signed(428, D_WIDTH),
        to_signed(434, D_WIDTH),
        to_signed(439, D_WIDTH),
        to_signed(445, D_WIDTH),
        to_signed(450, D_WIDTH),
        to_signed(455, D_WIDTH),
        to_signed(460, D_WIDTH),
        to_signed(464, D_WIDTH),
        to_signed(469, D_WIDTH),
        to_signed(474, D_WIDTH),
        to_signed(478, D_WIDTH),
        to_signed(482, D_WIDTH),
        to_signed(486, D_WIDTH),
        to_signed(490, D_WIDTH),
        to_signed(494, D_WIDTH),
        to_signed(498, D_WIDTH),
        to_signed(501, D_WIDTH),
        to_signed(504, D_WIDTH),
        to_signed(508, D_WIDTH),
        to_signed(511, D_WIDTH),
        to_signed(513, D_WIDTH),
        to_signed(516, D_WIDTH),
        to_signed(519, D_WIDTH),
        to_signed(521, D_WIDTH),
        to_signed(523, D_WIDTH),
        to_signed(525, D_WIDTH),
        to_signed(527, D_WIDTH),
        to_signed(529, D_WIDTH),
        to_signed(530, D_WIDTH),
        to_signed(531, D_WIDTH),
        to_signed(533, D_WIDTH),
        to_signed(533, D_WIDTH),
        to_signed(534, D_WIDTH),
        to_signed(535, D_WIDTH),
        to_signed(535, D_WIDTH),
        to_signed(535, D_WIDTH),
        to_signed(535, D_WIDTH),
        to_signed(535, D_WIDTH),
        to_signed(535, D_WIDTH),
        to_signed(534, D_WIDTH),
        to_signed(534, D_WIDTH),
        to_signed(533, D_WIDTH),
        to_signed(531, D_WIDTH),
        to_signed(530, D_WIDTH),
        to_signed(529, D_WIDTH),
        to_signed(527, D_WIDTH),
        to_signed(525, D_WIDTH),
        to_signed(523, D_WIDTH),
        to_signed(520, D_WIDTH),
        to_signed(518, D_WIDTH),
        to_signed(515, D_WIDTH),
        to_signed(512, D_WIDTH),
        to_signed(509, D_WIDTH),
        to_signed(506, D_WIDTH),
        to_signed(502, D_WIDTH),
        to_signed(498, D_WIDTH),
        to_signed(494, D_WIDTH),
        to_signed(490, D_WIDTH),
        to_signed(486, D_WIDTH),
        to_signed(481, D_WIDTH),
        to_signed(477, D_WIDTH),
        to_signed(472, D_WIDTH),
        to_signed(466, D_WIDTH),
        to_signed(461, D_WIDTH),
        to_signed(456, D_WIDTH),
        to_signed(450, D_WIDTH),
        to_signed(444, D_WIDTH),
        to_signed(438, D_WIDTH),
        to_signed(431, D_WIDTH),
        to_signed(425, D_WIDTH),
        to_signed(418, D_WIDTH),
        to_signed(411, D_WIDTH),
        to_signed(404, D_WIDTH),
        to_signed(397, D_WIDTH),
        to_signed(389, D_WIDTH),
        to_signed(382, D_WIDTH),
        to_signed(374, D_WIDTH),
        to_signed(366, D_WIDTH),
        to_signed(357, D_WIDTH),
        to_signed(349, D_WIDTH),
        to_signed(340, D_WIDTH),
        to_signed(332, D_WIDTH),
        to_signed(323, D_WIDTH),
        to_signed(314, D_WIDTH),
        to_signed(304, D_WIDTH),
        to_signed(295, D_WIDTH),
        to_signed(285, D_WIDTH),
        to_signed(275, D_WIDTH),
        to_signed(265, D_WIDTH),
        to_signed(255, D_WIDTH),
        to_signed(245, D_WIDTH),
        to_signed(235, D_WIDTH),
        to_signed(224, D_WIDTH),
        to_signed(213, D_WIDTH),
        to_signed(202, D_WIDTH),
        to_signed(191, D_WIDTH),
        to_signed(180, D_WIDTH),
        to_signed(169, D_WIDTH),
        to_signed(158, D_WIDTH),
        to_signed(146, D_WIDTH),
        to_signed(134, D_WIDTH),
        to_signed(123, D_WIDTH),
        to_signed(111, D_WIDTH),
        to_signed(99, D_WIDTH),
        to_signed(87, D_WIDTH),
        to_signed(74, D_WIDTH),
        to_signed(62, D_WIDTH),
        to_signed(49, D_WIDTH),
        to_signed(37, D_WIDTH),
        to_signed(24, D_WIDTH),
        to_signed(12, D_WIDTH),
        to_signed(-1, D_WIDTH),
        to_signed(-14, D_WIDTH),
        to_signed(-27, D_WIDTH),
        to_signed(-40, D_WIDTH),
        to_signed(-53, D_WIDTH),
        to_signed(-66, D_WIDTH),
        to_signed(-80, D_WIDTH),
        to_signed(-93, D_WIDTH),
        to_signed(-106, D_WIDTH),
        to_signed(-120, D_WIDTH),
        to_signed(-133, D_WIDTH),
        to_signed(-147, D_WIDTH),
        to_signed(-160, D_WIDTH),
        to_signed(-174, D_WIDTH),
        to_signed(-187, D_WIDTH),
        to_signed(-201, D_WIDTH),
        to_signed(-214, D_WIDTH),
        to_signed(-228, D_WIDTH),
        to_signed(-242, D_WIDTH),
        to_signed(-255, D_WIDTH),
        to_signed(-269, D_WIDTH),
        to_signed(-283, D_WIDTH),
        to_signed(-296, D_WIDTH),
        to_signed(-310, D_WIDTH),
        to_signed(-323, D_WIDTH),
        to_signed(-337, D_WIDTH),
        to_signed(-350, D_WIDTH),
        to_signed(-364, D_WIDTH),
        to_signed(-377, D_WIDTH),
        to_signed(-390, D_WIDTH),
        to_signed(-404, D_WIDTH),
        to_signed(-417, D_WIDTH),
        to_signed(-430, D_WIDTH),
        to_signed(-443, D_WIDTH),
        to_signed(-456, D_WIDTH),
        to_signed(-469, D_WIDTH),
        to_signed(-482, D_WIDTH),
        to_signed(-495, D_WIDTH),
        to_signed(-507, D_WIDTH),
        to_signed(-520, D_WIDTH),
        to_signed(-532, D_WIDTH),
        to_signed(-545, D_WIDTH),
        to_signed(-557, D_WIDTH),
        to_signed(-569, D_WIDTH),
        to_signed(-581, D_WIDTH),
        to_signed(-593, D_WIDTH),
        to_signed(-605, D_WIDTH),
        to_signed(-616, D_WIDTH),
        to_signed(-628, D_WIDTH),
        to_signed(-639, D_WIDTH),
        to_signed(-650, D_WIDTH),
        to_signed(-661, D_WIDTH),
        to_signed(-672, D_WIDTH),
        to_signed(-682, D_WIDTH),
        to_signed(-693, D_WIDTH),
        to_signed(-703, D_WIDTH),
        to_signed(-713, D_WIDTH),
        to_signed(-723, D_WIDTH),
        to_signed(-733, D_WIDTH),
        to_signed(-742, D_WIDTH),
        to_signed(-751, D_WIDTH),
        to_signed(-760, D_WIDTH),
        to_signed(-769, D_WIDTH),
        to_signed(-778, D_WIDTH),
        to_signed(-786, D_WIDTH),
        to_signed(-795, D_WIDTH),
        to_signed(-803, D_WIDTH),
        to_signed(-810, D_WIDTH),
        to_signed(-818, D_WIDTH),
        to_signed(-825, D_WIDTH),
        to_signed(-832, D_WIDTH),
        to_signed(-839, D_WIDTH),
        to_signed(-845, D_WIDTH),
        to_signed(-852, D_WIDTH),
        to_signed(-857, D_WIDTH),
        to_signed(-863, D_WIDTH),
        to_signed(-869, D_WIDTH),
        to_signed(-874, D_WIDTH),
        to_signed(-879, D_WIDTH),
        to_signed(-883, D_WIDTH),
        to_signed(-888, D_WIDTH),
        to_signed(-892, D_WIDTH),
        to_signed(-895, D_WIDTH),
        to_signed(-899, D_WIDTH),
        to_signed(-902, D_WIDTH),
        to_signed(-905, D_WIDTH),
        to_signed(-907, D_WIDTH),
        to_signed(-909, D_WIDTH),
        to_signed(-911, D_WIDTH),
        to_signed(-913, D_WIDTH),
        to_signed(-914, D_WIDTH),
        to_signed(-915, D_WIDTH),
        to_signed(-916, D_WIDTH),
        to_signed(-916, D_WIDTH),
        to_signed(-916, D_WIDTH),
        to_signed(-916, D_WIDTH),
        to_signed(-915, D_WIDTH),
        to_signed(-914, D_WIDTH),
        to_signed(-913, D_WIDTH),
        to_signed(-912, D_WIDTH),
        to_signed(-910, D_WIDTH),
        to_signed(-907, D_WIDTH),
        to_signed(-905, D_WIDTH),
        to_signed(-902, D_WIDTH),
        to_signed(-899, D_WIDTH),
        to_signed(-895, D_WIDTH),
        to_signed(-891, D_WIDTH),
        to_signed(-887, D_WIDTH),
        to_signed(-882, D_WIDTH),
        to_signed(-877, D_WIDTH),
        to_signed(-872, D_WIDTH),
        to_signed(-866, D_WIDTH),
        to_signed(-860, D_WIDTH),
        to_signed(-854, D_WIDTH),
        to_signed(-847, D_WIDTH),
        to_signed(-840, D_WIDTH),
        to_signed(-833, D_WIDTH),
        to_signed(-825, D_WIDTH),
        to_signed(-817, D_WIDTH),
        to_signed(-809, D_WIDTH),
        to_signed(-800, D_WIDTH),
        to_signed(-791, D_WIDTH),
        to_signed(-782, D_WIDTH),
        to_signed(-772, D_WIDTH),
        to_signed(-762, D_WIDTH),
        to_signed(-752, D_WIDTH),
        to_signed(-741, D_WIDTH),
        to_signed(-730, D_WIDTH),
        to_signed(-719, D_WIDTH),
        to_signed(-707, D_WIDTH),
        to_signed(-695, D_WIDTH),
        to_signed(-683, D_WIDTH),
        to_signed(-670, D_WIDTH),
        to_signed(-657, D_WIDTH),
        to_signed(-644, D_WIDTH),
        to_signed(-630, D_WIDTH),
        to_signed(-617, D_WIDTH),
        to_signed(-603, D_WIDTH),
        to_signed(-588, D_WIDTH),
        to_signed(-573, D_WIDTH),
        to_signed(-558, D_WIDTH),
        to_signed(-543, D_WIDTH),
        to_signed(-528, D_WIDTH),
        to_signed(-512, D_WIDTH),
        to_signed(-496, D_WIDTH),
        to_signed(-479, D_WIDTH),
        to_signed(-463, D_WIDTH),
        to_signed(-446, D_WIDTH),
        to_signed(-429, D_WIDTH),
        to_signed(-411, D_WIDTH),
        to_signed(-394, D_WIDTH),
        to_signed(-376, D_WIDTH),
        to_signed(-358, D_WIDTH),
        to_signed(-339, D_WIDTH),
        to_signed(-321, D_WIDTH),
        to_signed(-302, D_WIDTH),
        to_signed(-283, D_WIDTH),
        to_signed(-264, D_WIDTH),
        to_signed(-244, D_WIDTH),
        to_signed(-225, D_WIDTH),
        to_signed(-205, D_WIDTH),
        to_signed(-185, D_WIDTH),
        to_signed(-165, D_WIDTH),
        to_signed(-144, D_WIDTH),
        to_signed(-124, D_WIDTH),
        to_signed(-103, D_WIDTH),
        to_signed(-82, D_WIDTH),
        to_signed(-61, D_WIDTH),
        to_signed(-40, D_WIDTH),
        to_signed(-19, D_WIDTH),
        to_signed(3, D_WIDTH),
        to_signed(24, D_WIDTH),
        to_signed(46, D_WIDTH),
        to_signed(67, D_WIDTH),
        to_signed(89, D_WIDTH),
        to_signed(111, D_WIDTH),
        to_signed(133, D_WIDTH),
        to_signed(155, D_WIDTH),
        to_signed(177, D_WIDTH),
        to_signed(200, D_WIDTH),
        to_signed(222, D_WIDTH),
        to_signed(244, D_WIDTH),
        to_signed(267, D_WIDTH),
        to_signed(289, D_WIDTH),
        to_signed(312, D_WIDTH),
        to_signed(334, D_WIDTH),
        to_signed(356, D_WIDTH),
        to_signed(379, D_WIDTH),
        to_signed(401, D_WIDTH),
        to_signed(424, D_WIDTH),
        to_signed(446, D_WIDTH),
        to_signed(469, D_WIDTH),
        to_signed(491, D_WIDTH),
        to_signed(513, D_WIDTH),
        to_signed(536, D_WIDTH),
        to_signed(558, D_WIDTH),
        to_signed(580, D_WIDTH),
        to_signed(602, D_WIDTH),
        to_signed(624, D_WIDTH),
        to_signed(646, D_WIDTH),
        to_signed(667, D_WIDTH),
        to_signed(689, D_WIDTH),
        to_signed(711, D_WIDTH),
        to_signed(732, D_WIDTH),
        to_signed(753, D_WIDTH),
        to_signed(774, D_WIDTH),
        to_signed(795, D_WIDTH),
        to_signed(816, D_WIDTH),
        to_signed(837, D_WIDTH),
        to_signed(857, D_WIDTH),
        to_signed(877, D_WIDTH),
        to_signed(897, D_WIDTH),
        to_signed(917, D_WIDTH),
        to_signed(937, D_WIDTH),
        to_signed(956, D_WIDTH),
        to_signed(975, D_WIDTH),
        to_signed(994, D_WIDTH),
        to_signed(1013, D_WIDTH),
        to_signed(1032, D_WIDTH),
        to_signed(1050, D_WIDTH),
        to_signed(1068, D_WIDTH),
        to_signed(1085, D_WIDTH),
        to_signed(1103, D_WIDTH),
        to_signed(1120, D_WIDTH),
        to_signed(1137, D_WIDTH),
        to_signed(1153, D_WIDTH),
        to_signed(1169, D_WIDTH),
        to_signed(1185, D_WIDTH),
        to_signed(1201, D_WIDTH),
        to_signed(1216, D_WIDTH),
        to_signed(1231, D_WIDTH),
        to_signed(1245, D_WIDTH),
        to_signed(1259, D_WIDTH),
        to_signed(1273, D_WIDTH),
        to_signed(1286, D_WIDTH),
        to_signed(1299, D_WIDTH),
        to_signed(1312, D_WIDTH),
        to_signed(1324, D_WIDTH),
        to_signed(1336, D_WIDTH),
        to_signed(1347, D_WIDTH),
        to_signed(1358, D_WIDTH),
        to_signed(1369, D_WIDTH),
        to_signed(1379, D_WIDTH),
        to_signed(1389, D_WIDTH),
        to_signed(1398, D_WIDTH),
        to_signed(1407, D_WIDTH),
        to_signed(1415, D_WIDTH),
        to_signed(1423, D_WIDTH),
        to_signed(1431, D_WIDTH),
        to_signed(1438, D_WIDTH),
        to_signed(1445, D_WIDTH),
        to_signed(1451, D_WIDTH),
        to_signed(1456, D_WIDTH),
        to_signed(1461, D_WIDTH),
        to_signed(1466, D_WIDTH),
        to_signed(1470, D_WIDTH),
        to_signed(1474, D_WIDTH),
        to_signed(1477, D_WIDTH),
        to_signed(1480, D_WIDTH),
        to_signed(1482, D_WIDTH),
        to_signed(1484, D_WIDTH),
        to_signed(1485, D_WIDTH),
        to_signed(1486, D_WIDTH),
        to_signed(1486, D_WIDTH),
        to_signed(1485, D_WIDTH),
        to_signed(1484, D_WIDTH),
        to_signed(1483, D_WIDTH),
        to_signed(1481, D_WIDTH),
        to_signed(1478, D_WIDTH),
        to_signed(1475, D_WIDTH),
        to_signed(1472, D_WIDTH),
        to_signed(1468, D_WIDTH),
        to_signed(1463, D_WIDTH),
        to_signed(1458, D_WIDTH),
        to_signed(1452, D_WIDTH),
        to_signed(1446, D_WIDTH),
        to_signed(1439, D_WIDTH),
        to_signed(1432, D_WIDTH),
        to_signed(1424, D_WIDTH),
        to_signed(1415, D_WIDTH),
        to_signed(1406, D_WIDTH),
        to_signed(1397, D_WIDTH),
        to_signed(1387, D_WIDTH),
        to_signed(1376, D_WIDTH),
        to_signed(1365, D_WIDTH),
        to_signed(1354, D_WIDTH),
        to_signed(1341, D_WIDTH),
        to_signed(1329, D_WIDTH),
        to_signed(1315, D_WIDTH),
        to_signed(1301, D_WIDTH),
        to_signed(1287, D_WIDTH),
        to_signed(1272, D_WIDTH),
        to_signed(1257, D_WIDTH),
        to_signed(1241, D_WIDTH),
        to_signed(1225, D_WIDTH),
        to_signed(1208, D_WIDTH),
        to_signed(1190, D_WIDTH),
        to_signed(1172, D_WIDTH),
        to_signed(1154, D_WIDTH),
        to_signed(1135, D_WIDTH),
        to_signed(1115, D_WIDTH),
        to_signed(1095, D_WIDTH),
        to_signed(1075, D_WIDTH),
        to_signed(1054, D_WIDTH),
        to_signed(1032, D_WIDTH),
        to_signed(1010, D_WIDTH),
        to_signed(988, D_WIDTH),
        to_signed(965, D_WIDTH),
        to_signed(942, D_WIDTH),
        to_signed(918, D_WIDTH),
        to_signed(894, D_WIDTH),
        to_signed(869, D_WIDTH),
        to_signed(844, D_WIDTH),
        to_signed(819, D_WIDTH),
        to_signed(793, D_WIDTH),
        to_signed(766, D_WIDTH),
        to_signed(740, D_WIDTH),
        to_signed(712, D_WIDTH),
        to_signed(685, D_WIDTH),
        to_signed(657, D_WIDTH),
        to_signed(629, D_WIDTH),
        to_signed(600, D_WIDTH),
        to_signed(571, D_WIDTH),
        to_signed(542, D_WIDTH),
        to_signed(512, D_WIDTH),
        to_signed(482, D_WIDTH),
        to_signed(451, D_WIDTH),
        to_signed(421, D_WIDTH),
        to_signed(390, D_WIDTH),
        to_signed(358, D_WIDTH),
        to_signed(327, D_WIDTH),
        to_signed(295, D_WIDTH),
        to_signed(263, D_WIDTH),
        to_signed(230, D_WIDTH),
        to_signed(197, D_WIDTH),
        to_signed(165, D_WIDTH),
        to_signed(131, D_WIDTH),
        to_signed(98, D_WIDTH),
        to_signed(64, D_WIDTH),
        to_signed(31, D_WIDTH),
        to_signed(-3, D_WIDTH),
        to_signed(-37, D_WIDTH),
        to_signed(-72, D_WIDTH),
        to_signed(-106, D_WIDTH),
        to_signed(-141, D_WIDTH),
        to_signed(-175, D_WIDTH),
        to_signed(-210, D_WIDTH),
        to_signed(-245, D_WIDTH),
        to_signed(-280, D_WIDTH),
        to_signed(-315, D_WIDTH),
        to_signed(-351, D_WIDTH),
        to_signed(-386, D_WIDTH),
        to_signed(-421, D_WIDTH),
        to_signed(-457, D_WIDTH),
        to_signed(-492, D_WIDTH),
        to_signed(-527, D_WIDTH),
        to_signed(-563, D_WIDTH),
        to_signed(-598, D_WIDTH),
        to_signed(-633, D_WIDTH),
        to_signed(-669, D_WIDTH),
        to_signed(-704, D_WIDTH),
        to_signed(-739, D_WIDTH),
        to_signed(-774, D_WIDTH),
        to_signed(-809, D_WIDTH),
        to_signed(-844, D_WIDTH),
        to_signed(-879, D_WIDTH),
        to_signed(-914, D_WIDTH),
        to_signed(-948, D_WIDTH),
        to_signed(-983, D_WIDTH),
        to_signed(-1017, D_WIDTH),
        to_signed(-1051, D_WIDTH),
        to_signed(-1085, D_WIDTH),
        to_signed(-1118, D_WIDTH),
        to_signed(-1152, D_WIDTH),
        to_signed(-1185, D_WIDTH),
        to_signed(-1218, D_WIDTH),
        to_signed(-1250, D_WIDTH),
        to_signed(-1283, D_WIDTH),
        to_signed(-1315, D_WIDTH),
        to_signed(-1347, D_WIDTH),
        to_signed(-1378, D_WIDTH),
        to_signed(-1410, D_WIDTH),
        to_signed(-1440, D_WIDTH),
        to_signed(-1471, D_WIDTH),
        to_signed(-1501, D_WIDTH),
        to_signed(-1531, D_WIDTH),
        to_signed(-1560, D_WIDTH),
        to_signed(-1589, D_WIDTH),
        to_signed(-1618, D_WIDTH),
        to_signed(-1646, D_WIDTH),
        to_signed(-1674, D_WIDTH),
        to_signed(-1701, D_WIDTH),
        to_signed(-1728, D_WIDTH),
        to_signed(-1754, D_WIDTH),
        to_signed(-1780, D_WIDTH),
        to_signed(-1806, D_WIDTH),
        to_signed(-1831, D_WIDTH),
        to_signed(-1855, D_WIDTH),
        to_signed(-1879, D_WIDTH),
        to_signed(-1902, D_WIDTH),
        to_signed(-1925, D_WIDTH),
        to_signed(-1947, D_WIDTH),
        to_signed(-1969, D_WIDTH),
        to_signed(-1990, D_WIDTH),
        to_signed(-2011, D_WIDTH),
        to_signed(-2030, D_WIDTH),
        to_signed(-2050, D_WIDTH),
        to_signed(-2068, D_WIDTH),
        to_signed(-2087, D_WIDTH),
        to_signed(-2104, D_WIDTH),
        to_signed(-2121, D_WIDTH),
        to_signed(-2137, D_WIDTH),
        to_signed(-2152, D_WIDTH),
        to_signed(-2167, D_WIDTH),
        to_signed(-2181, D_WIDTH),
        to_signed(-2195, D_WIDTH),
        to_signed(-2207, D_WIDTH),
        to_signed(-2219, D_WIDTH),
        to_signed(-2230, D_WIDTH),
        to_signed(-2241, D_WIDTH),
        to_signed(-2251, D_WIDTH),
        to_signed(-2260, D_WIDTH),
        to_signed(-2268, D_WIDTH),
        to_signed(-2276, D_WIDTH),
        to_signed(-2283, D_WIDTH),
        to_signed(-2289, D_WIDTH),
        to_signed(-2294, D_WIDTH),
        to_signed(-2299, D_WIDTH),
        to_signed(-2302, D_WIDTH),
        to_signed(-2305, D_WIDTH),
        to_signed(-2307, D_WIDTH),
        to_signed(-2309, D_WIDTH),
        to_signed(-2309, D_WIDTH),
        to_signed(-2309, D_WIDTH),
        to_signed(-2308, D_WIDTH),
        to_signed(-2306, D_WIDTH),
        to_signed(-2304, D_WIDTH),
        to_signed(-2300, D_WIDTH),
        to_signed(-2296, D_WIDTH),
        to_signed(-2291, D_WIDTH),
        to_signed(-2285, D_WIDTH),
        to_signed(-2278, D_WIDTH),
        to_signed(-2270, D_WIDTH),
        to_signed(-2262, D_WIDTH),
        to_signed(-2253, D_WIDTH),
        to_signed(-2243, D_WIDTH),
        to_signed(-2232, D_WIDTH),
        to_signed(-2220, D_WIDTH),
        to_signed(-2207, D_WIDTH),
        to_signed(-2194, D_WIDTH),
        to_signed(-2180, D_WIDTH),
        to_signed(-2165, D_WIDTH),
        to_signed(-2149, D_WIDTH),
        to_signed(-2132, D_WIDTH),
        to_signed(-2114, D_WIDTH),
        to_signed(-2096, D_WIDTH),
        to_signed(-2077, D_WIDTH),
        to_signed(-2057, D_WIDTH),
        to_signed(-2036, D_WIDTH),
        to_signed(-2014, D_WIDTH),
        to_signed(-1991, D_WIDTH),
        to_signed(-1968, D_WIDTH),
        to_signed(-1944, D_WIDTH),
        to_signed(-1919, D_WIDTH),
        to_signed(-1893, D_WIDTH),
        to_signed(-1867, D_WIDTH),
        to_signed(-1840, D_WIDTH),
        to_signed(-1812, D_WIDTH),
        to_signed(-1783, D_WIDTH),
        to_signed(-1753, D_WIDTH),
        to_signed(-1723, D_WIDTH),
        to_signed(-1692, D_WIDTH),
        to_signed(-1660, D_WIDTH),
        to_signed(-1627, D_WIDTH),
        to_signed(-1594, D_WIDTH),
        to_signed(-1560, D_WIDTH),
        to_signed(-1525, D_WIDTH),
        to_signed(-1490, D_WIDTH),
        to_signed(-1454, D_WIDTH),
        to_signed(-1417, D_WIDTH),
        to_signed(-1379, D_WIDTH),
        to_signed(-1341, D_WIDTH),
        to_signed(-1302, D_WIDTH),
        to_signed(-1263, D_WIDTH),
        to_signed(-1223, D_WIDTH),
        to_signed(-1182, D_WIDTH),
        to_signed(-1141, D_WIDTH),
        to_signed(-1099, D_WIDTH),
        to_signed(-1056, D_WIDTH),
        to_signed(-1013, D_WIDTH),
        to_signed(-969, D_WIDTH),
        to_signed(-925, D_WIDTH),
        to_signed(-880, D_WIDTH),
        to_signed(-835, D_WIDTH),
        to_signed(-789, D_WIDTH),
        to_signed(-743, D_WIDTH),
        to_signed(-696, D_WIDTH),
        to_signed(-649, D_WIDTH),
        to_signed(-601, D_WIDTH),
        to_signed(-553, D_WIDTH),
        to_signed(-504, D_WIDTH),
        to_signed(-455, D_WIDTH),
        to_signed(-406, D_WIDTH),
        to_signed(-356, D_WIDTH),
        to_signed(-306, D_WIDTH),
        to_signed(-255, D_WIDTH),
        to_signed(-204, D_WIDTH),
        to_signed(-153, D_WIDTH),
        to_signed(-102, D_WIDTH),
        to_signed(-50, D_WIDTH),
        to_signed(2, D_WIDTH),
        to_signed(55, D_WIDTH),
        to_signed(107, D_WIDTH),
        to_signed(160, D_WIDTH),
        to_signed(213, D_WIDTH),
        to_signed(266, D_WIDTH),
        to_signed(319, D_WIDTH),
        to_signed(373, D_WIDTH),
        to_signed(427, D_WIDTH),
        to_signed(480, D_WIDTH),
        to_signed(534, D_WIDTH),
        to_signed(588, D_WIDTH),
        to_signed(642, D_WIDTH),
        to_signed(696, D_WIDTH),
        to_signed(750, D_WIDTH),
        to_signed(804, D_WIDTH),
        to_signed(858, D_WIDTH),
        to_signed(912, D_WIDTH),
        to_signed(966, D_WIDTH),
        to_signed(1020, D_WIDTH),
        to_signed(1074, D_WIDTH),
        to_signed(1127, D_WIDTH),
        to_signed(1181, D_WIDTH),
        to_signed(1234, D_WIDTH),
        to_signed(1287, D_WIDTH),
        to_signed(1340, D_WIDTH),
        to_signed(1393, D_WIDTH),
        to_signed(1446, D_WIDTH),
        to_signed(1498, D_WIDTH),
        to_signed(1550, D_WIDTH),
        to_signed(1602, D_WIDTH),
        to_signed(1654, D_WIDTH),
        to_signed(1705, D_WIDTH),
        to_signed(1756, D_WIDTH),
        to_signed(1806, D_WIDTH),
        to_signed(1856, D_WIDTH),
        to_signed(1906, D_WIDTH),
        to_signed(1955, D_WIDTH),
        to_signed(2004, D_WIDTH),
        to_signed(2052, D_WIDTH),
        to_signed(2100, D_WIDTH),
        to_signed(2147, D_WIDTH),
        to_signed(2194, D_WIDTH),
        to_signed(2241, D_WIDTH),
        to_signed(2286, D_WIDTH),
        to_signed(2332, D_WIDTH),
        to_signed(2376, D_WIDTH),
        to_signed(2420, D_WIDTH),
        to_signed(2463, D_WIDTH),
        to_signed(2506, D_WIDTH),
        to_signed(2548, D_WIDTH),
        to_signed(2590, D_WIDTH),
        to_signed(2630, D_WIDTH),
        to_signed(2670, D_WIDTH),
        to_signed(2709, D_WIDTH),
        to_signed(2748, D_WIDTH),
        to_signed(2786, D_WIDTH),
        to_signed(2823, D_WIDTH),
        to_signed(2859, D_WIDTH),
        to_signed(2894, D_WIDTH),
        to_signed(2928, D_WIDTH),
        to_signed(2962, D_WIDTH),
        to_signed(2995, D_WIDTH),
        to_signed(3027, D_WIDTH),
        to_signed(3058, D_WIDTH),
        to_signed(3088, D_WIDTH),
        to_signed(3117, D_WIDTH),
        to_signed(3145, D_WIDTH),
        to_signed(3172, D_WIDTH),
        to_signed(3198, D_WIDTH),
        to_signed(3224, D_WIDTH),
        to_signed(3248, D_WIDTH),
        to_signed(3271, D_WIDTH),
        to_signed(3293, D_WIDTH),
        to_signed(3314, D_WIDTH),
        to_signed(3335, D_WIDTH),
        to_signed(3354, D_WIDTH),
        to_signed(3372, D_WIDTH),
        to_signed(3389, D_WIDTH),
        to_signed(3404, D_WIDTH),
        to_signed(3419, D_WIDTH),
        to_signed(3433, D_WIDTH),
        to_signed(3445, D_WIDTH),
        to_signed(3456, D_WIDTH),
        to_signed(3467, D_WIDTH),
        to_signed(3476, D_WIDTH),
        to_signed(3483, D_WIDTH),
        to_signed(3490, D_WIDTH),
        to_signed(3496, D_WIDTH),
        to_signed(3500, D_WIDTH),
        to_signed(3503, D_WIDTH),
        to_signed(3505, D_WIDTH),
        to_signed(3506, D_WIDTH),
        to_signed(3505, D_WIDTH),
        to_signed(3503, D_WIDTH),
        to_signed(3500, D_WIDTH),
        to_signed(3496, D_WIDTH),
        to_signed(3491, D_WIDTH),
        to_signed(3484, D_WIDTH),
        to_signed(3476, D_WIDTH),
        to_signed(3467, D_WIDTH),
        to_signed(3456, D_WIDTH),
        to_signed(3445, D_WIDTH),
        to_signed(3432, D_WIDTH),
        to_signed(3418, D_WIDTH),
        to_signed(3402, D_WIDTH),
        to_signed(3385, D_WIDTH),
        to_signed(3368, D_WIDTH),
        to_signed(3348, D_WIDTH),
        to_signed(3328, D_WIDTH),
        to_signed(3306, D_WIDTH),
        to_signed(3283, D_WIDTH),
        to_signed(3259, D_WIDTH),
        to_signed(3233, D_WIDTH),
        to_signed(3207, D_WIDTH),
        to_signed(3179, D_WIDTH),
        to_signed(3149, D_WIDTH),
        to_signed(3119, D_WIDTH),
        to_signed(3087, D_WIDTH),
        to_signed(3054, D_WIDTH),
        to_signed(3020, D_WIDTH),
        to_signed(2985, D_WIDTH),
        to_signed(2948, D_WIDTH),
        to_signed(2910, D_WIDTH),
        to_signed(2871, D_WIDTH),
        to_signed(2831, D_WIDTH),
        to_signed(2790, D_WIDTH),
        to_signed(2747, D_WIDTH),
        to_signed(2704, D_WIDTH),
        to_signed(2659, D_WIDTH),
        to_signed(2613, D_WIDTH),
        to_signed(2566, D_WIDTH),
        to_signed(2517, D_WIDTH),
        to_signed(2468, D_WIDTH),
        to_signed(2418, D_WIDTH),
        to_signed(2366, D_WIDTH),
        to_signed(2313, D_WIDTH),
        to_signed(2260, D_WIDTH),
        to_signed(2205, D_WIDTH),
        to_signed(2149, D_WIDTH),
        to_signed(2093, D_WIDTH),
        to_signed(2035, D_WIDTH),
        to_signed(1976, D_WIDTH),
        to_signed(1916, D_WIDTH),
        to_signed(1856, D_WIDTH),
        to_signed(1794, D_WIDTH),
        to_signed(1731, D_WIDTH),
        to_signed(1668, D_WIDTH),
        to_signed(1604, D_WIDTH),
        to_signed(1538, D_WIDTH),
        to_signed(1472, D_WIDTH),
        to_signed(1405, D_WIDTH),
        to_signed(1338, D_WIDTH),
        to_signed(1269, D_WIDTH),
        to_signed(1200, D_WIDTH),
        to_signed(1130, D_WIDTH),
        to_signed(1059, D_WIDTH),
        to_signed(987, D_WIDTH),
        to_signed(915, D_WIDTH),
        to_signed(842, D_WIDTH),
        to_signed(769, D_WIDTH),
        to_signed(695, D_WIDTH),
        to_signed(620, D_WIDTH),
        to_signed(545, D_WIDTH),
        to_signed(469, D_WIDTH),
        to_signed(392, D_WIDTH),
        to_signed(315, D_WIDTH),
        to_signed(238, D_WIDTH),
        to_signed(160, D_WIDTH),
        to_signed(82, D_WIDTH),
        to_signed(3, D_WIDTH),
        to_signed(-76, D_WIDTH),
        to_signed(-156, D_WIDTH),
        to_signed(-235, D_WIDTH),
        to_signed(-316, D_WIDTH),
        to_signed(-396, D_WIDTH),
        to_signed(-477, D_WIDTH),
        to_signed(-558, D_WIDTH),
        to_signed(-639, D_WIDTH),
        to_signed(-720, D_WIDTH),
        to_signed(-801, D_WIDTH),
        to_signed(-883, D_WIDTH),
        to_signed(-965, D_WIDTH),
        to_signed(-1046, D_WIDTH),
        to_signed(-1128, D_WIDTH),
        to_signed(-1210, D_WIDTH),
        to_signed(-1292, D_WIDTH),
        to_signed(-1373, D_WIDTH),
        to_signed(-1455, D_WIDTH),
        to_signed(-1536, D_WIDTH),
        to_signed(-1618, D_WIDTH),
        to_signed(-1699, D_WIDTH),
        to_signed(-1780, D_WIDTH),
        to_signed(-1861, D_WIDTH),
        to_signed(-1941, D_WIDTH),
        to_signed(-2022, D_WIDTH),
        to_signed(-2102, D_WIDTH),
        to_signed(-2181, D_WIDTH),
        to_signed(-2261, D_WIDTH),
        to_signed(-2339, D_WIDTH),
        to_signed(-2418, D_WIDTH),
        to_signed(-2496, D_WIDTH),
        to_signed(-2573, D_WIDTH),
        to_signed(-2650, D_WIDTH),
        to_signed(-2727, D_WIDTH),
        to_signed(-2803, D_WIDTH),
        to_signed(-2878, D_WIDTH),
        to_signed(-2953, D_WIDTH),
        to_signed(-3027, D_WIDTH),
        to_signed(-3100, D_WIDTH),
        to_signed(-3173, D_WIDTH),
        to_signed(-3245, D_WIDTH),
        to_signed(-3316, D_WIDTH),
        to_signed(-3386, D_WIDTH),
        to_signed(-3456, D_WIDTH),
        to_signed(-3524, D_WIDTH),
        to_signed(-3592, D_WIDTH),
        to_signed(-3659, D_WIDTH),
        to_signed(-3725, D_WIDTH),
        to_signed(-3790, D_WIDTH),
        to_signed(-3854, D_WIDTH),
        to_signed(-3917, D_WIDTH),
        to_signed(-3978, D_WIDTH),
        to_signed(-4039, D_WIDTH),
        to_signed(-4099, D_WIDTH),
        to_signed(-4158, D_WIDTH),
        to_signed(-4215, D_WIDTH),
        to_signed(-4271, D_WIDTH),
        to_signed(-4326, D_WIDTH),
        to_signed(-4380, D_WIDTH),
        to_signed(-4433, D_WIDTH),
        to_signed(-4484, D_WIDTH),
        to_signed(-4534, D_WIDTH),
        to_signed(-4583, D_WIDTH),
        to_signed(-4630, D_WIDTH),
        to_signed(-4676, D_WIDTH),
        to_signed(-4720, D_WIDTH),
        to_signed(-4764, D_WIDTH),
        to_signed(-4805, D_WIDTH),
        to_signed(-4846, D_WIDTH),
        to_signed(-4884, D_WIDTH),
        to_signed(-4922, D_WIDTH),
        to_signed(-4957, D_WIDTH),
        to_signed(-4992, D_WIDTH),
        to_signed(-5024, D_WIDTH),
        to_signed(-5055, D_WIDTH),
        to_signed(-5085, D_WIDTH),
        to_signed(-5112, D_WIDTH),
        to_signed(-5139, D_WIDTH),
        to_signed(-5163, D_WIDTH),
        to_signed(-5186, D_WIDTH),
        to_signed(-5207, D_WIDTH),
        to_signed(-5227, D_WIDTH),
        to_signed(-5245, D_WIDTH),
        to_signed(-5261, D_WIDTH),
        to_signed(-5275, D_WIDTH),
        to_signed(-5288, D_WIDTH),
        to_signed(-5298, D_WIDTH),
        to_signed(-5307, D_WIDTH),
        to_signed(-5315, D_WIDTH),
        to_signed(-5320, D_WIDTH),
        to_signed(-5323, D_WIDTH),
        to_signed(-5325, D_WIDTH),
        to_signed(-5325, D_WIDTH),
        to_signed(-5323, D_WIDTH),
        to_signed(-5319, D_WIDTH),
        to_signed(-5314, D_WIDTH),
        to_signed(-5306, D_WIDTH),
        to_signed(-5297, D_WIDTH),
        to_signed(-5285, D_WIDTH),
        to_signed(-5272, D_WIDTH),
        to_signed(-5257, D_WIDTH),
        to_signed(-5240, D_WIDTH),
        to_signed(-5221, D_WIDTH),
        to_signed(-5200, D_WIDTH),
        to_signed(-5178, D_WIDTH),
        to_signed(-5153, D_WIDTH),
        to_signed(-5127, D_WIDTH),
        to_signed(-5098, D_WIDTH),
        to_signed(-5068, D_WIDTH),
        to_signed(-5035, D_WIDTH),
        to_signed(-5001, D_WIDTH),
        to_signed(-4965, D_WIDTH),
        to_signed(-4927, D_WIDTH),
        to_signed(-4887, D_WIDTH),
        to_signed(-4845, D_WIDTH),
        to_signed(-4802, D_WIDTH),
        to_signed(-4756, D_WIDTH),
        to_signed(-4708, D_WIDTH),
        to_signed(-4659, D_WIDTH),
        to_signed(-4608, D_WIDTH),
        to_signed(-4555, D_WIDTH),
        to_signed(-4500, D_WIDTH),
        to_signed(-4443, D_WIDTH),
        to_signed(-4384, D_WIDTH),
        to_signed(-4324, D_WIDTH),
        to_signed(-4262, D_WIDTH),
        to_signed(-4198, D_WIDTH),
        to_signed(-4132, D_WIDTH),
        to_signed(-4064, D_WIDTH),
        to_signed(-3995, D_WIDTH),
        to_signed(-3924, D_WIDTH),
        to_signed(-3851, D_WIDTH),
        to_signed(-3776, D_WIDTH),
        to_signed(-3700, D_WIDTH),
        to_signed(-3622, D_WIDTH),
        to_signed(-3542, D_WIDTH),
        to_signed(-3461, D_WIDTH),
        to_signed(-3378, D_WIDTH),
        to_signed(-3294, D_WIDTH),
        to_signed(-3208, D_WIDTH),
        to_signed(-3120, D_WIDTH),
        to_signed(-3031, D_WIDTH),
        to_signed(-2940, D_WIDTH),
        to_signed(-2848, D_WIDTH),
        to_signed(-2754, D_WIDTH),
        to_signed(-2659, D_WIDTH),
        to_signed(-2563, D_WIDTH),
        to_signed(-2465, D_WIDTH),
        to_signed(-2365, D_WIDTH),
        to_signed(-2265, D_WIDTH),
        to_signed(-2163, D_WIDTH),
        to_signed(-2059, D_WIDTH),
        to_signed(-1955, D_WIDTH),
        to_signed(-1849, D_WIDTH),
        to_signed(-1742, D_WIDTH),
        to_signed(-1634, D_WIDTH),
        to_signed(-1525, D_WIDTH),
        to_signed(-1415, D_WIDTH),
        to_signed(-1303, D_WIDTH),
        to_signed(-1191, D_WIDTH),
        to_signed(-1077, D_WIDTH),
        to_signed(-963, D_WIDTH),
        to_signed(-848, D_WIDTH),
        to_signed(-731, D_WIDTH),
        to_signed(-614, D_WIDTH),
        to_signed(-496, D_WIDTH),
        to_signed(-377, D_WIDTH),
        to_signed(-258, D_WIDTH),
        to_signed(-138, D_WIDTH),
        to_signed(-17, D_WIDTH),
        to_signed(105, D_WIDTH),
        to_signed(227, D_WIDTH),
        to_signed(350, D_WIDTH),
        to_signed(473, D_WIDTH),
        to_signed(597, D_WIDTH),
        to_signed(722, D_WIDTH),
        to_signed(846, D_WIDTH),
        to_signed(971, D_WIDTH),
        to_signed(1097, D_WIDTH),
        to_signed(1223, D_WIDTH),
        to_signed(1349, D_WIDTH),
        to_signed(1475, D_WIDTH),
        to_signed(1601, D_WIDTH),
        to_signed(1728, D_WIDTH),
        to_signed(1854, D_WIDTH),
        to_signed(1981, D_WIDTH),
        to_signed(2108, D_WIDTH),
        to_signed(2234, D_WIDTH),
        to_signed(2361, D_WIDTH),
        to_signed(2487, D_WIDTH),
        to_signed(2613, D_WIDTH),
        to_signed(2739, D_WIDTH),
        to_signed(2865, D_WIDTH),
        to_signed(2990, D_WIDTH),
        to_signed(3115, D_WIDTH),
        to_signed(3240, D_WIDTH),
        to_signed(3364, D_WIDTH),
        to_signed(3488, D_WIDTH),
        to_signed(3611, D_WIDTH),
        to_signed(3734, D_WIDTH),
        to_signed(3856, D_WIDTH),
        to_signed(3977, D_WIDTH),
        to_signed(4098, D_WIDTH),
        to_signed(4218, D_WIDTH),
        to_signed(4337, D_WIDTH),
        to_signed(4455, D_WIDTH),
        to_signed(4572, D_WIDTH),
        to_signed(4689, D_WIDTH),
        to_signed(4804, D_WIDTH),
        to_signed(4919, D_WIDTH),
        to_signed(5032, D_WIDTH),
        to_signed(5144, D_WIDTH),
        to_signed(5255, D_WIDTH),
        to_signed(5365, D_WIDTH),
        to_signed(5474, D_WIDTH),
        to_signed(5581, D_WIDTH),
        to_signed(5687, D_WIDTH),
        to_signed(5792, D_WIDTH),
        to_signed(5895, D_WIDTH),
        to_signed(5997, D_WIDTH),
        to_signed(6097, D_WIDTH),
        to_signed(6196, D_WIDTH),
        to_signed(6293, D_WIDTH),
        to_signed(6388, D_WIDTH),
        to_signed(6482, D_WIDTH),
        to_signed(6574, D_WIDTH),
        to_signed(6664, D_WIDTH),
        to_signed(6753, D_WIDTH),
        to_signed(6839, D_WIDTH),
        to_signed(6924, D_WIDTH),
        to_signed(7007, D_WIDTH),
        to_signed(7088, D_WIDTH),
        to_signed(7167, D_WIDTH),
        to_signed(7244, D_WIDTH),
        to_signed(7319, D_WIDTH),
        to_signed(7391, D_WIDTH),
        to_signed(7462, D_WIDTH),
        to_signed(7530, D_WIDTH),
        to_signed(7596, D_WIDTH),
        to_signed(7660, D_WIDTH),
        to_signed(7722, D_WIDTH),
        to_signed(7781, D_WIDTH),
        to_signed(7838, D_WIDTH),
        to_signed(7893, D_WIDTH),
        to_signed(7945, D_WIDTH),
        to_signed(7995, D_WIDTH),
        to_signed(8042, D_WIDTH),
        to_signed(8087, D_WIDTH),
        to_signed(8129, D_WIDTH),
        to_signed(8168, D_WIDTH),
        to_signed(8205, D_WIDTH),
        to_signed(8240, D_WIDTH),
        to_signed(8271, D_WIDTH),
        to_signed(8300, D_WIDTH),
        to_signed(8327, D_WIDTH),
        to_signed(8350, D_WIDTH),
        to_signed(8371, D_WIDTH),
        to_signed(8389, D_WIDTH),
        to_signed(8404, D_WIDTH),
        to_signed(8417, D_WIDTH),
        to_signed(8427, D_WIDTH),
        to_signed(8433, D_WIDTH),
        to_signed(8437, D_WIDTH),
        to_signed(8438, D_WIDTH),
        to_signed(8436, D_WIDTH),
        to_signed(8431, D_WIDTH),
        to_signed(8423, D_WIDTH),
        to_signed(8412, D_WIDTH),
        to_signed(8399, D_WIDTH),
        to_signed(8382, D_WIDTH),
        to_signed(8362, D_WIDTH),
        to_signed(8339, D_WIDTH),
        to_signed(8313, D_WIDTH),
        to_signed(8284, D_WIDTH),
        to_signed(8252, D_WIDTH),
        to_signed(8217, D_WIDTH),
        to_signed(8179, D_WIDTH),
        to_signed(8138, D_WIDTH),
        to_signed(8094, D_WIDTH),
        to_signed(8047, D_WIDTH),
        to_signed(7997, D_WIDTH),
        to_signed(7943, D_WIDTH),
        to_signed(7887, D_WIDTH),
        to_signed(7827, D_WIDTH),
        to_signed(7764, D_WIDTH),
        to_signed(7699, D_WIDTH),
        to_signed(7630, D_WIDTH),
        to_signed(7558, D_WIDTH),
        to_signed(7483, D_WIDTH),
        to_signed(7405, D_WIDTH),
        to_signed(7324, D_WIDTH),
        to_signed(7240, D_WIDTH),
        to_signed(7153, D_WIDTH),
        to_signed(7063, D_WIDTH),
        to_signed(6970, D_WIDTH),
        to_signed(6873, D_WIDTH),
        to_signed(6774, D_WIDTH),
        to_signed(6672, D_WIDTH),
        to_signed(6567, D_WIDTH),
        to_signed(6459, D_WIDTH),
        to_signed(6348, D_WIDTH),
        to_signed(6234, D_WIDTH),
        to_signed(6118, D_WIDTH),
        to_signed(5998, D_WIDTH),
        to_signed(5876, D_WIDTH),
        to_signed(5750, D_WIDTH),
        to_signed(5622, D_WIDTH),
        to_signed(5492, D_WIDTH),
        to_signed(5358, D_WIDTH),
        to_signed(5222, D_WIDTH),
        to_signed(5083, D_WIDTH),
        to_signed(4942, D_WIDTH),
        to_signed(4797, D_WIDTH),
        to_signed(4651, D_WIDTH),
        to_signed(4501, D_WIDTH),
        to_signed(4349, D_WIDTH),
        to_signed(4195, D_WIDTH),
        to_signed(4038, D_WIDTH),
        to_signed(3879, D_WIDTH),
        to_signed(3717, D_WIDTH),
        to_signed(3553, D_WIDTH),
        to_signed(3387, D_WIDTH),
        to_signed(3219, D_WIDTH),
        to_signed(3048, D_WIDTH),
        to_signed(2875, D_WIDTH),
        to_signed(2700, D_WIDTH),
        to_signed(2523, D_WIDTH),
        to_signed(2343, D_WIDTH),
        to_signed(2162, D_WIDTH),
        to_signed(1979, D_WIDTH),
        to_signed(1794, D_WIDTH),
        to_signed(1607, D_WIDTH),
        to_signed(1418, D_WIDTH),
        to_signed(1227, D_WIDTH),
        to_signed(1035, D_WIDTH),
        to_signed(841, D_WIDTH),
        to_signed(646, D_WIDTH),
        to_signed(449, D_WIDTH),
        to_signed(250, D_WIDTH),
        to_signed(50, D_WIDTH),
        to_signed(-151, D_WIDTH),
        to_signed(-354, D_WIDTH),
        to_signed(-558, D_WIDTH),
        to_signed(-763, D_WIDTH),
        to_signed(-969, D_WIDTH),
        to_signed(-1177, D_WIDTH),
        to_signed(-1385, D_WIDTH),
        to_signed(-1594, D_WIDTH),
        to_signed(-1805, D_WIDTH),
        to_signed(-2016, D_WIDTH),
        to_signed(-2228, D_WIDTH),
        to_signed(-2440, D_WIDTH),
        to_signed(-2654, D_WIDTH),
        to_signed(-2867, D_WIDTH),
        to_signed(-3082, D_WIDTH),
        to_signed(-3296, D_WIDTH),
        to_signed(-3512, D_WIDTH),
        to_signed(-3727, D_WIDTH),
        to_signed(-3943, D_WIDTH),
        to_signed(-4159, D_WIDTH),
        to_signed(-4374, D_WIDTH),
        to_signed(-4590, D_WIDTH),
        to_signed(-4806, D_WIDTH),
        to_signed(-5022, D_WIDTH),
        to_signed(-5238, D_WIDTH),
        to_signed(-5453, D_WIDTH),
        to_signed(-5668, D_WIDTH),
        to_signed(-5883, D_WIDTH),
        to_signed(-6097, D_WIDTH),
        to_signed(-6311, D_WIDTH),
        to_signed(-6524, D_WIDTH),
        to_signed(-6736, D_WIDTH),
        to_signed(-6947, D_WIDTH),
        to_signed(-7158, D_WIDTH),
        to_signed(-7368, D_WIDTH),
        to_signed(-7576, D_WIDTH),
        to_signed(-7784, D_WIDTH),
        to_signed(-7991, D_WIDTH),
        to_signed(-8196, D_WIDTH),
        to_signed(-8400, D_WIDTH),
        to_signed(-8602, D_WIDTH),
        to_signed(-8804, D_WIDTH),
        to_signed(-9003, D_WIDTH),
        to_signed(-9201, D_WIDTH),
        to_signed(-9397, D_WIDTH),
        to_signed(-9592, D_WIDTH),
        to_signed(-9785, D_WIDTH),
        to_signed(-9975, D_WIDTH),
        to_signed(-10164, D_WIDTH),
        to_signed(-10351, D_WIDTH),
        to_signed(-10535, D_WIDTH),
        to_signed(-10717, D_WIDTH),
        to_signed(-10897, D_WIDTH),
        to_signed(-11075, D_WIDTH),
        to_signed(-11250, D_WIDTH),
        to_signed(-11423, D_WIDTH),
        to_signed(-11593, D_WIDTH),
        to_signed(-11760, D_WIDTH),
        to_signed(-11925, D_WIDTH),
        to_signed(-12087, D_WIDTH),
        to_signed(-12245, D_WIDTH),
        to_signed(-12401, D_WIDTH),
        to_signed(-12554, D_WIDTH),
        to_signed(-12704, D_WIDTH),
        to_signed(-12850, D_WIDTH),
        to_signed(-12993, D_WIDTH),
        to_signed(-13133, D_WIDTH),
        to_signed(-13269, D_WIDTH),
        to_signed(-13402, D_WIDTH),
        to_signed(-13532, D_WIDTH),
        to_signed(-13657, D_WIDTH),
        to_signed(-13779, D_WIDTH),
        to_signed(-13898, D_WIDTH),
        to_signed(-14012, D_WIDTH),
        to_signed(-14123, D_WIDTH),
        to_signed(-14229, D_WIDTH),
        to_signed(-14331, D_WIDTH),
        to_signed(-14430, D_WIDTH),
        to_signed(-14524, D_WIDTH),
        to_signed(-14614, D_WIDTH),
        to_signed(-14699, D_WIDTH),
        to_signed(-14781, D_WIDTH),
        to_signed(-14857, D_WIDTH),
        to_signed(-14930, D_WIDTH),
        to_signed(-14997, D_WIDTH),
        to_signed(-15061, D_WIDTH),
        to_signed(-15119, D_WIDTH),
        to_signed(-15173, D_WIDTH),
        to_signed(-15222, D_WIDTH),
        to_signed(-15266, D_WIDTH),
        to_signed(-15305, D_WIDTH),
        to_signed(-15339, D_WIDTH),
        to_signed(-15368, D_WIDTH),
        to_signed(-15392, D_WIDTH),
        to_signed(-15411, D_WIDTH),
        to_signed(-15425, D_WIDTH),
        to_signed(-15433, D_WIDTH),
        to_signed(-15437, D_WIDTH),
        to_signed(-15435, D_WIDTH),
        to_signed(-15427, D_WIDTH),
        to_signed(-15414, D_WIDTH),
        to_signed(-15396, D_WIDTH),
        to_signed(-15372, D_WIDTH),
        to_signed(-15343, D_WIDTH),
        to_signed(-15308, D_WIDTH),
        to_signed(-15267, D_WIDTH),
        to_signed(-15221, D_WIDTH),
        to_signed(-15169, D_WIDTH),
        to_signed(-15112, D_WIDTH),
        to_signed(-15048, D_WIDTH),
        to_signed(-14979, D_WIDTH),
        to_signed(-14904, D_WIDTH),
        to_signed(-14823, D_WIDTH),
        to_signed(-14736, D_WIDTH),
        to_signed(-14643, D_WIDTH),
        to_signed(-14544, D_WIDTH),
        to_signed(-14440, D_WIDTH),
        to_signed(-14329, D_WIDTH),
        to_signed(-14212, D_WIDTH),
        to_signed(-14089, D_WIDTH),
        to_signed(-13960, D_WIDTH),
        to_signed(-13825, D_WIDTH),
        to_signed(-13684, D_WIDTH),
        to_signed(-13537, D_WIDTH),
        to_signed(-13383, D_WIDTH),
        to_signed(-13224, D_WIDTH),
        to_signed(-13058, D_WIDTH),
        to_signed(-12886, D_WIDTH),
        to_signed(-12708, D_WIDTH),
        to_signed(-12523, D_WIDTH),
        to_signed(-12333, D_WIDTH),
        to_signed(-12136, D_WIDTH),
        to_signed(-11933, D_WIDTH),
        to_signed(-11724, D_WIDTH),
        to_signed(-11508, D_WIDTH),
        to_signed(-11287, D_WIDTH),
        to_signed(-11059, D_WIDTH),
        to_signed(-10825, D_WIDTH),
        to_signed(-10585, D_WIDTH),
        to_signed(-10338, D_WIDTH),
        to_signed(-10085, D_WIDTH),
        to_signed(-9827, D_WIDTH),
        to_signed(-9562, D_WIDTH),
        to_signed(-9290, D_WIDTH),
        to_signed(-9013, D_WIDTH),
        to_signed(-8730, D_WIDTH),
        to_signed(-8440, D_WIDTH),
        to_signed(-8144, D_WIDTH),
        to_signed(-7843, D_WIDTH),
        to_signed(-7535, D_WIDTH),
        to_signed(-7221, D_WIDTH),
        to_signed(-6901, D_WIDTH),
        to_signed(-6576, D_WIDTH),
        to_signed(-6244, D_WIDTH),
        to_signed(-5906, D_WIDTH),
        to_signed(-5563, D_WIDTH),
        to_signed(-5214, D_WIDTH),
        to_signed(-4858, D_WIDTH),
        to_signed(-4498, D_WIDTH),
        to_signed(-4131, D_WIDTH),
        to_signed(-3759, D_WIDTH),
        to_signed(-3381, D_WIDTH),
        to_signed(-2997, D_WIDTH),
        to_signed(-2608, D_WIDTH),
        to_signed(-2213, D_WIDTH),
        to_signed(-1813, D_WIDTH),
        to_signed(-1407, D_WIDTH),
        to_signed(-996, D_WIDTH),
        to_signed(-580, D_WIDTH),
        to_signed(-159, D_WIDTH),
        to_signed(268, D_WIDTH),
        to_signed(700, D_WIDTH),
        to_signed(1137, D_WIDTH),
        to_signed(1580, D_WIDTH),
        to_signed(2027, D_WIDTH),
        to_signed(2479, D_WIDTH),
        to_signed(2936, D_WIDTH),
        to_signed(3397, D_WIDTH),
        to_signed(3864, D_WIDTH),
        to_signed(4335, D_WIDTH),
        to_signed(4811, D_WIDTH),
        to_signed(5291, D_WIDTH),
        to_signed(5776, D_WIDTH),
        to_signed(6265, D_WIDTH),
        to_signed(6759, D_WIDTH),
        to_signed(7256, D_WIDTH),
        to_signed(7758, D_WIDTH),
        to_signed(8264, D_WIDTH),
        to_signed(8774, D_WIDTH),
        to_signed(9288, D_WIDTH),
        to_signed(9806, D_WIDTH),
        to_signed(10328, D_WIDTH),
        to_signed(10853, D_WIDTH),
        to_signed(11382, D_WIDTH),
        to_signed(11914, D_WIDTH),
        to_signed(12450, D_WIDTH),
        to_signed(12989, D_WIDTH),
        to_signed(13532, D_WIDTH),
        to_signed(14078, D_WIDTH),
        to_signed(14626, D_WIDTH),
        to_signed(15178, D_WIDTH),
        to_signed(15733, D_WIDTH),
        to_signed(16290, D_WIDTH),
        to_signed(16850, D_WIDTH),
        to_signed(17413, D_WIDTH),
        to_signed(17978, D_WIDTH),
        to_signed(18546, D_WIDTH),
        to_signed(19116, D_WIDTH),
        to_signed(19688, D_WIDTH),
        to_signed(20263, D_WIDTH),
        to_signed(20839, D_WIDTH),
        to_signed(21417, D_WIDTH),
        to_signed(21998, D_WIDTH),
        to_signed(22579, D_WIDTH),
        to_signed(23163, D_WIDTH),
        to_signed(23748, D_WIDTH),
        to_signed(24334, D_WIDTH),
        to_signed(24922, D_WIDTH),
        to_signed(25511, D_WIDTH),
        to_signed(26101, D_WIDTH),
        to_signed(26692, D_WIDTH),
        to_signed(27284, D_WIDTH),
        to_signed(27877, D_WIDTH),
        to_signed(28470, D_WIDTH),
        to_signed(29064, D_WIDTH),
        to_signed(29658, D_WIDTH),
        to_signed(30253, D_WIDTH),
        to_signed(30848, D_WIDTH),
        to_signed(31443, D_WIDTH),
        to_signed(32038, D_WIDTH),
        to_signed(32632, D_WIDTH),
        to_signed(33227, D_WIDTH),
        to_signed(33821, D_WIDTH),
        to_signed(34415, D_WIDTH),
        to_signed(35008, D_WIDTH),
        to_signed(35601, D_WIDTH),
        to_signed(36193, D_WIDTH),
        to_signed(36784, D_WIDTH),
        to_signed(37374, D_WIDTH),
        to_signed(37963, D_WIDTH),
        to_signed(38550, D_WIDTH),
        to_signed(39137, D_WIDTH),
        to_signed(39721, D_WIDTH),
        to_signed(40305, D_WIDTH),
        to_signed(40886, D_WIDTH),
        to_signed(41466, D_WIDTH),
        to_signed(42044, D_WIDTH),
        to_signed(42619, D_WIDTH),
        to_signed(43193, D_WIDTH),
        to_signed(43764, D_WIDTH),
        to_signed(44334, D_WIDTH),
        to_signed(44900, D_WIDTH),
        to_signed(45464, D_WIDTH),
        to_signed(46025, D_WIDTH),
        to_signed(46584, D_WIDTH),
        to_signed(47139, D_WIDTH),
        to_signed(47692, D_WIDTH),
        to_signed(48241, D_WIDTH),
        to_signed(48788, D_WIDTH),
        to_signed(49330, D_WIDTH),
        to_signed(49870, D_WIDTH),
        to_signed(50406, D_WIDTH),
        to_signed(50938, D_WIDTH),
        to_signed(51466, D_WIDTH),
        to_signed(51991, D_WIDTH),
        to_signed(52511, D_WIDTH),
        to_signed(53027, D_WIDTH),
        to_signed(53540, D_WIDTH),
        to_signed(54048, D_WIDTH),
        to_signed(54551, D_WIDTH),
        to_signed(55050, D_WIDTH),
        to_signed(55544, D_WIDTH),
        to_signed(56034, D_WIDTH),
        to_signed(56519, D_WIDTH),
        to_signed(56999, D_WIDTH),
        to_signed(57474, D_WIDTH),
        to_signed(57944, D_WIDTH),
        to_signed(58408, D_WIDTH),
        to_signed(58868, D_WIDTH),
        to_signed(59322, D_WIDTH),
        to_signed(59770, D_WIDTH),
        to_signed(60213, D_WIDTH),
        to_signed(60650, D_WIDTH),
        to_signed(61082, D_WIDTH),
        to_signed(61508, D_WIDTH),
        to_signed(61927, D_WIDTH),
        to_signed(62341, D_WIDTH),
        to_signed(62749, D_WIDTH),
        to_signed(63150, D_WIDTH),
        to_signed(63546, D_WIDTH),
        to_signed(63934, D_WIDTH),
        to_signed(64317, D_WIDTH),
        to_signed(64693, D_WIDTH),
        to_signed(65062, D_WIDTH),
        to_signed(65425, D_WIDTH),
        to_signed(65781, D_WIDTH),
        to_signed(66130, D_WIDTH),
        to_signed(66473, D_WIDTH),
        to_signed(66808, D_WIDTH),
        to_signed(67136, D_WIDTH),
        to_signed(67458, D_WIDTH),
        to_signed(67772, D_WIDTH),
        to_signed(68079, D_WIDTH),
        to_signed(68378, D_WIDTH),
        to_signed(68671, D_WIDTH),
        to_signed(68955, D_WIDTH),
        to_signed(69233, D_WIDTH),
        to_signed(69503, D_WIDTH),
        to_signed(69765, D_WIDTH),
        to_signed(70020, D_WIDTH),
        to_signed(70267, D_WIDTH),
        to_signed(70506, D_WIDTH),
        to_signed(70738, D_WIDTH),
        to_signed(70961, D_WIDTH),
        to_signed(71177, D_WIDTH),
        to_signed(71385, D_WIDTH),
        to_signed(71585, D_WIDTH),
        to_signed(71777, D_WIDTH),
        to_signed(71961, D_WIDTH),
        to_signed(72136, D_WIDTH),
        to_signed(72304, D_WIDTH),
        to_signed(72463, D_WIDTH),
        to_signed(72615, D_WIDTH),
        to_signed(72758, D_WIDTH),
        to_signed(72892, D_WIDTH),
        to_signed(73019, D_WIDTH),
        to_signed(73137, D_WIDTH),
        to_signed(73247, D_WIDTH),
        to_signed(73348, D_WIDTH),
        to_signed(73441, D_WIDTH),
        to_signed(73526, D_WIDTH),
        to_signed(73602, D_WIDTH),
        to_signed(73670, D_WIDTH),
        to_signed(73730, D_WIDTH),
        to_signed(73781, D_WIDTH),
        to_signed(73823, D_WIDTH),
        to_signed(73857, D_WIDTH),
        to_signed(73882, D_WIDTH),
        to_signed(73899, D_WIDTH),
        to_signed(73908, D_WIDTH),
        -- 2048 - 1920 = 128 padding works
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH),
        to_signed(0, D_WIDTH)
    );

begin

    process(clk)
    begin
        if rising_edge(clk) then
            if clk_en = '1' then
                data <= coeff_list(to_integer(addr));
            end if;
        end if;
    end process;

end rtl;
